magic
tech sky130B
magscale 1 2
timestamp 1667873852
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 137830 700816 137836 700868
rect 137888 700856 137894 700868
rect 157334 700856 157340 700868
rect 137888 700828 157340 700856
rect 137888 700816 137894 700828
rect 157334 700816 157340 700828
rect 157392 700816 157398 700868
rect 155954 700748 155960 700800
rect 156012 700788 156018 700800
rect 202782 700788 202788 700800
rect 156012 700760 202788 700788
rect 156012 700748 156018 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 160738 700720 160744 700732
rect 89220 700692 160744 700720
rect 89220 700680 89226 700692
rect 160738 700680 160744 700692
rect 160796 700680 160802 700732
rect 154574 700612 154580 700664
rect 154632 700652 154638 700664
rect 267642 700652 267648 700664
rect 154632 700624 267648 700652
rect 154632 700612 154638 700624
rect 267642 700612 267648 700624
rect 267700 700612 267706 700664
rect 24302 700544 24308 700596
rect 24360 700584 24366 700596
rect 162210 700584 162216 700596
rect 24360 700556 162216 700584
rect 24360 700544 24366 700556
rect 162210 700544 162216 700556
rect 162268 700544 162274 700596
rect 8110 700476 8116 700528
rect 8168 700516 8174 700528
rect 162118 700516 162124 700528
rect 8168 700488 162124 700516
rect 8168 700476 8174 700488
rect 162118 700476 162124 700488
rect 162176 700476 162182 700528
rect 153286 700408 153292 700460
rect 153344 700448 153350 700460
rect 332502 700448 332508 700460
rect 153344 700420 332508 700448
rect 153344 700408 153350 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 152458 700340 152464 700392
rect 152516 700380 152522 700392
rect 413646 700380 413652 700392
rect 152516 700352 413652 700380
rect 152516 700340 152522 700352
rect 413646 700340 413652 700352
rect 413704 700340 413710 700392
rect 489178 700340 489184 700392
rect 489236 700380 489242 700392
rect 527174 700380 527180 700392
rect 489236 700352 527180 700380
rect 489236 700340 489242 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 527818 700340 527824 700392
rect 527876 700380 527882 700392
rect 559650 700380 559656 700392
rect 527876 700352 559656 700380
rect 527876 700340 527882 700352
rect 559650 700340 559656 700352
rect 559708 700340 559714 700392
rect 148318 700272 148324 700324
rect 148376 700312 148382 700324
rect 543458 700312 543464 700324
rect 148376 700284 543464 700312
rect 148376 700272 148382 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 396718 699660 396724 699712
rect 396776 699700 396782 699712
rect 397454 699700 397460 699712
rect 396776 699672 397460 699700
rect 396776 699660 396782 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 428458 699660 428464 699712
rect 428516 699700 428522 699712
rect 429838 699700 429844 699712
rect 428516 699672 429844 699700
rect 428516 699660 428522 699672
rect 429838 699660 429844 699672
rect 429896 699660 429902 699712
rect 146294 696940 146300 696992
rect 146352 696980 146358 696992
rect 580166 696980 580172 696992
rect 146352 696952 580172 696980
rect 146352 696940 146358 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683204 3424 683256
rect 3476 683244 3482 683256
rect 161474 683244 161480 683256
rect 3476 683216 161480 683244
rect 3476 683204 3482 683216
rect 161474 683204 161480 683216
rect 161532 683204 161538 683256
rect 146938 683136 146944 683188
rect 146996 683176 147002 683188
rect 580166 683176 580172 683188
rect 146996 683148 580172 683176
rect 146996 683136 147002 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 163498 670732 163504 670744
rect 3568 670704 163504 670732
rect 3568 670692 3574 670704
rect 163498 670692 163504 670704
rect 163556 670692 163562 670744
rect 498838 670692 498844 670744
rect 498896 670732 498902 670744
rect 580166 670732 580172 670744
rect 498896 670704 580172 670732
rect 498896 670692 498902 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 163590 656928 163596 656940
rect 3476 656900 163596 656928
rect 3476 656888 3482 656900
rect 163590 656888 163596 656900
rect 163648 656888 163654 656940
rect 182818 643084 182824 643136
rect 182876 643124 182882 643136
rect 580166 643124 580172 643136
rect 182876 643096 580172 643124
rect 182876 643084 182882 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 164234 632108 164240 632120
rect 3476 632080 164240 632108
rect 3476 632068 3482 632080
rect 164234 632068 164240 632080
rect 164292 632068 164298 632120
rect 188338 630640 188344 630692
rect 188396 630680 188402 630692
rect 580166 630680 580172 630692
rect 188396 630652 580172 630680
rect 188396 630640 188402 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 164878 618304 164884 618316
rect 3200 618276 164884 618304
rect 3200 618264 3206 618276
rect 164878 618264 164884 618276
rect 164936 618264 164942 618316
rect 143626 616836 143632 616888
rect 143684 616876 143690 616888
rect 580166 616876 580172 616888
rect 143684 616848 580172 616876
rect 143684 616836 143690 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 164970 605860 164976 605872
rect 3292 605832 164976 605860
rect 3292 605820 3298 605832
rect 164970 605820 164976 605832
rect 165028 605820 165034 605872
rect 142430 590656 142436 590708
rect 142488 590696 142494 590708
rect 579798 590696 579804 590708
rect 142488 590668 579804 590696
rect 142488 590656 142494 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 165614 579680 165620 579692
rect 3384 579652 165620 579680
rect 3384 579640 3390 579652
rect 165614 579640 165620 579652
rect 165672 579640 165678 579692
rect 144178 576852 144184 576904
rect 144236 576892 144242 576904
rect 580166 576892 580172 576904
rect 144236 576864 580172 576892
rect 144236 576852 144242 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 167638 565876 167644 565888
rect 3476 565848 167644 565876
rect 3476 565836 3482 565848
rect 167638 565836 167644 565848
rect 167696 565836 167702 565888
rect 142798 563048 142804 563100
rect 142856 563088 142862 563100
rect 579798 563088 579804 563100
rect 142856 563060 579804 563088
rect 142856 563048 142862 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 166258 553432 166264 553444
rect 3476 553404 166264 553432
rect 3476 553392 3482 553404
rect 166258 553392 166264 553404
rect 166316 553392 166322 553444
rect 181438 536800 181444 536852
rect 181496 536840 181502 536852
rect 580166 536840 580172 536852
rect 181496 536812 580172 536840
rect 181496 536800 181502 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 166994 527184 167000 527196
rect 3476 527156 167000 527184
rect 3476 527144 3482 527156
rect 166994 527144 167000 527156
rect 167052 527144 167058 527196
rect 142890 524424 142896 524476
rect 142948 524464 142954 524476
rect 580166 524464 580172 524476
rect 142948 524436 580172 524464
rect 142948 524424 142954 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 7558 514808 7564 514820
rect 3476 514780 7564 514808
rect 3476 514768 3482 514780
rect 7558 514768 7564 514780
rect 7616 514768 7622 514820
rect 180058 510620 180064 510672
rect 180116 510660 180122 510672
rect 580166 510660 580172 510672
rect 180116 510632 580172 510660
rect 180116 510620 180122 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 167730 501004 167736 501016
rect 3108 500976 167736 501004
rect 3108 500964 3114 500976
rect 167730 500964 167736 500976
rect 167788 500964 167794 501016
rect 139578 484372 139584 484424
rect 139636 484412 139642 484424
rect 580166 484412 580172 484424
rect 139636 484384 580172 484412
rect 139636 484372 139642 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 140038 470568 140044 470620
rect 140096 470608 140102 470620
rect 579982 470608 579988 470620
rect 140096 470580 579988 470608
rect 140096 470568 140102 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 170398 462380 170404 462392
rect 3568 462352 170404 462380
rect 3568 462340 3574 462352
rect 170398 462340 170404 462352
rect 170456 462340 170462 462392
rect 178678 456764 178684 456816
rect 178736 456804 178742 456816
rect 580166 456804 580172 456816
rect 178736 456776 580172 456804
rect 178736 456764 178742 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 157426 450508 157432 450560
rect 157484 450548 157490 450560
rect 169754 450548 169760 450560
rect 157484 450520 169760 450548
rect 157484 450508 157490 450520
rect 169754 450508 169760 450520
rect 169812 450508 169818 450560
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 170490 448576 170496 448588
rect 3200 448548 170496 448576
rect 3200 448536 3206 448548
rect 170490 448536 170496 448548
rect 170548 448536 170554 448588
rect 138658 430584 138664 430636
rect 138716 430624 138722 430636
rect 580166 430624 580172 430636
rect 138716 430596 580172 430624
rect 138716 430584 138722 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 169754 422328 169760 422340
rect 3568 422300 169760 422328
rect 3568 422288 3574 422300
rect 169754 422288 169760 422300
rect 169812 422288 169818 422340
rect 138750 418140 138756 418192
rect 138808 418180 138814 418192
rect 580166 418180 580172 418192
rect 138808 418152 580172 418180
rect 138808 418140 138814 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 171778 409884 171784 409896
rect 2924 409856 171784 409884
rect 2924 409844 2930 409856
rect 171778 409844 171784 409856
rect 171836 409844 171842 409896
rect 185578 404336 185584 404388
rect 185636 404376 185642 404388
rect 580166 404376 580172 404388
rect 185636 404348 580172 404376
rect 185636 404336 185642 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 171870 397508 171876 397520
rect 3568 397480 171876 397508
rect 3568 397468 3574 397480
rect 171870 397468 171876 397480
rect 171928 397468 171934 397520
rect 196618 378156 196624 378208
rect 196676 378196 196682 378208
rect 580166 378196 580172 378208
rect 196676 378168 580172 378196
rect 196676 378156 196682 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 2774 371288 2780 371340
rect 2832 371328 2838 371340
rect 4798 371328 4804 371340
rect 2832 371300 4804 371328
rect 2832 371288 2838 371300
rect 4798 371288 4804 371300
rect 4856 371288 4862 371340
rect 3510 358368 3516 358420
rect 3568 358408 3574 358420
rect 8938 358408 8944 358420
rect 3568 358380 8944 358408
rect 3568 358368 3574 358380
rect 8938 358368 8944 358380
rect 8996 358368 9002 358420
rect 135254 351908 135260 351960
rect 135312 351948 135318 351960
rect 580166 351948 580172 351960
rect 135312 351920 580172 351948
rect 135312 351908 135318 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 149698 345080 149704 345092
rect 3384 345052 149704 345080
rect 3384 345040 3390 345052
rect 149698 345040 149704 345052
rect 149756 345040 149762 345092
rect 134518 324300 134524 324352
rect 134576 324340 134582 324352
rect 580166 324340 580172 324352
rect 134576 324312 580172 324340
rect 134576 324300 134582 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3326 318792 3332 318844
rect 3384 318832 3390 318844
rect 173894 318832 173900 318844
rect 3384 318804 173900 318832
rect 3384 318792 3390 318804
rect 173894 318792 173900 318804
rect 173952 318792 173958 318844
rect 135898 311856 135904 311908
rect 135956 311896 135962 311908
rect 579982 311896 579988 311908
rect 135956 311868 579988 311896
rect 135956 311856 135962 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 3510 304988 3516 305040
rect 3568 305028 3574 305040
rect 175918 305028 175924 305040
rect 3568 305000 175924 305028
rect 3568 304988 3574 305000
rect 175918 304988 175924 305000
rect 175976 304988 175982 305040
rect 134610 298120 134616 298172
rect 134668 298160 134674 298172
rect 580166 298160 580172 298172
rect 134668 298132 580172 298160
rect 134668 298120 134674 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 174538 292584 174544 292596
rect 3568 292556 174544 292584
rect 3568 292544 3574 292556
rect 174538 292544 174544 292556
rect 174596 292544 174602 292596
rect 145558 289076 145564 289128
rect 145616 289116 145622 289128
rect 188338 289116 188344 289128
rect 145616 289088 188344 289116
rect 145616 289076 145622 289088
rect 188338 289076 188344 289088
rect 188396 289076 188402 289128
rect 149054 287648 149060 287700
rect 149112 287688 149118 287700
rect 462314 287688 462320 287700
rect 149112 287660 462320 287688
rect 149112 287648 149118 287660
rect 462314 287648 462320 287660
rect 462372 287648 462378 287700
rect 137278 286288 137284 286340
rect 137336 286328 137342 286340
rect 196618 286328 196624 286340
rect 137336 286300 196624 286328
rect 137336 286288 137342 286300
rect 196618 286288 196624 286300
rect 196676 286288 196682 286340
rect 150434 284928 150440 284980
rect 150492 284968 150498 284980
rect 396718 284968 396724 284980
rect 150492 284940 396724 284968
rect 150492 284928 150498 284940
rect 396718 284928 396724 284940
rect 396776 284928 396782 284980
rect 189442 283568 189448 283620
rect 189500 283608 189506 283620
rect 489178 283608 489184 283620
rect 189500 283580 489184 283608
rect 189500 283568 189506 283580
rect 489178 283568 489184 283580
rect 489236 283568 489242 283620
rect 147674 282888 147680 282940
rect 147732 282928 147738 282940
rect 189074 282928 189080 282940
rect 147732 282900 189080 282928
rect 147732 282888 147738 282900
rect 189074 282888 189080 282900
rect 189132 282928 189138 282940
rect 189442 282928 189448 282940
rect 189132 282900 189448 282928
rect 189132 282888 189138 282900
rect 189442 282888 189448 282900
rect 189500 282888 189506 282940
rect 144914 282140 144920 282192
rect 144972 282180 144978 282192
rect 182818 282180 182824 282192
rect 144972 282152 182824 282180
rect 144972 282140 144978 282152
rect 182818 282140 182824 282152
rect 182876 282140 182882 282192
rect 140774 280780 140780 280832
rect 140832 280820 140838 280832
rect 181438 280820 181444 280832
rect 140832 280792 181444 280820
rect 140832 280780 140838 280792
rect 181438 280780 181444 280792
rect 181496 280780 181502 280832
rect 40034 279420 40040 279472
rect 40092 279460 40098 279472
rect 160094 279460 160100 279472
rect 40092 279432 160100 279460
rect 40092 279420 40098 279432
rect 160094 279420 160100 279432
rect 160152 279420 160158 279472
rect 151078 275272 151084 275324
rect 151136 275312 151142 275324
rect 428458 275312 428464 275324
rect 151136 275284 428464 275312
rect 151136 275272 151142 275284
rect 428458 275272 428464 275284
rect 428516 275272 428522 275324
rect 8938 273912 8944 273964
rect 8996 273952 9002 273964
rect 173158 273952 173164 273964
rect 8996 273924 173164 273952
rect 8996 273912 9002 273924
rect 173158 273912 173164 273924
rect 173216 273912 173222 273964
rect 187694 273912 187700 273964
rect 187752 273952 187758 273964
rect 364334 273952 364340 273964
rect 187752 273924 364340 273952
rect 187752 273912 187758 273924
rect 364334 273912 364340 273924
rect 364392 273912 364398 273964
rect 151814 273232 151820 273284
rect 151872 273272 151878 273284
rect 187694 273272 187700 273284
rect 151872 273244 187700 273272
rect 151872 273232 151878 273244
rect 187694 273232 187700 273244
rect 187752 273232 187758 273284
rect 133138 271872 133144 271924
rect 133196 271912 133202 271924
rect 580166 271912 580172 271924
rect 133196 271884 580172 271912
rect 133196 271872 133202 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 7558 271192 7564 271244
rect 7616 271232 7622 271244
rect 169018 271232 169024 271244
rect 7616 271204 169024 271232
rect 7616 271192 7622 271204
rect 169018 271192 169024 271204
rect 169076 271192 169082 271244
rect 149146 271124 149152 271176
rect 149204 271164 149210 271176
rect 494054 271164 494060 271176
rect 149204 271136 494060 271164
rect 149204 271124 149210 271136
rect 494054 271124 494060 271136
rect 494112 271124 494118 271176
rect 71774 269832 71780 269884
rect 71832 269872 71838 269884
rect 158806 269872 158812 269884
rect 71832 269844 158812 269872
rect 71832 269832 71838 269844
rect 158806 269832 158812 269844
rect 158864 269832 158870 269884
rect 147766 269764 147772 269816
rect 147824 269804 147830 269816
rect 527818 269804 527824 269816
rect 147824 269776 527824 269804
rect 147824 269764 147830 269776
rect 527818 269764 527824 269776
rect 527876 269764 527882 269816
rect 4798 268404 4804 268456
rect 4856 268444 4862 268456
rect 172514 268444 172520 268456
rect 4856 268416 172520 268444
rect 4856 268404 4862 268416
rect 172514 268404 172520 268416
rect 172572 268404 172578 268456
rect 146202 268336 146208 268388
rect 146260 268376 146266 268388
rect 498838 268376 498844 268388
rect 146260 268348 498844 268376
rect 146260 268336 146266 268348
rect 498838 268336 498844 268348
rect 498896 268336 498902 268388
rect 137830 266976 137836 267028
rect 137888 267016 137894 267028
rect 185578 267016 185584 267028
rect 137888 266988 185584 267016
rect 137888 266976 137894 266988
rect 185578 266976 185584 266988
rect 185636 266976 185642 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 175918 266404 175924 266416
rect 3108 266376 175924 266404
rect 3108 266364 3114 266376
rect 175918 266364 175924 266376
rect 175976 266364 175982 266416
rect 141418 265684 141424 265736
rect 141476 265724 141482 265736
rect 180058 265724 180064 265736
rect 141476 265696 180064 265724
rect 141476 265684 141482 265696
rect 180058 265684 180064 265696
rect 180116 265684 180122 265736
rect 3418 265616 3424 265668
rect 3476 265656 3482 265668
rect 169202 265656 169208 265668
rect 3476 265628 169208 265656
rect 3476 265616 3482 265628
rect 169202 265616 169208 265628
rect 169260 265616 169266 265668
rect 172514 265548 172520 265600
rect 172572 265588 172578 265600
rect 190454 265588 190460 265600
rect 172572 265560 190460 265588
rect 172572 265548 172578 265560
rect 190454 265548 190460 265560
rect 190512 265548 190518 265600
rect 171870 265480 171876 265532
rect 171928 265520 171934 265532
rect 190822 265520 190828 265532
rect 171928 265492 190828 265520
rect 171928 265480 171934 265492
rect 190822 265480 190828 265492
rect 190880 265480 190886 265532
rect 174538 265412 174544 265464
rect 174596 265452 174602 265464
rect 194870 265452 194876 265464
rect 174596 265424 194876 265452
rect 174596 265412 174602 265424
rect 194870 265412 194876 265424
rect 194928 265412 194934 265464
rect 175826 265344 175832 265396
rect 175884 265384 175890 265396
rect 196434 265384 196440 265396
rect 175884 265356 196440 265384
rect 175884 265344 175890 265356
rect 196434 265344 196440 265356
rect 196492 265344 196498 265396
rect 170214 265276 170220 265328
rect 170272 265316 170278 265328
rect 170490 265316 170496 265328
rect 170272 265288 170496 265316
rect 170272 265276 170278 265288
rect 170490 265276 170496 265288
rect 170548 265316 170554 265328
rect 192018 265316 192024 265328
rect 170548 265288 192024 265316
rect 170548 265276 170554 265288
rect 192018 265276 192024 265288
rect 192076 265276 192082 265328
rect 171686 265208 171692 265260
rect 171744 265248 171750 265260
rect 171870 265248 171876 265260
rect 171744 265220 171876 265248
rect 171744 265208 171750 265220
rect 171870 265208 171876 265220
rect 171928 265208 171934 265260
rect 173342 265208 173348 265260
rect 173400 265248 173406 265260
rect 197630 265248 197636 265260
rect 173400 265220 197636 265248
rect 173400 265208 173406 265220
rect 197630 265208 197636 265220
rect 197688 265208 197694 265260
rect 171778 265140 171784 265192
rect 171836 265180 171842 265192
rect 196526 265180 196532 265192
rect 171836 265152 196532 265180
rect 171836 265140 171842 265152
rect 196526 265140 196532 265152
rect 196584 265140 196590 265192
rect 169110 265072 169116 265124
rect 169168 265112 169174 265124
rect 196250 265112 196256 265124
rect 169168 265084 196256 265112
rect 169168 265072 169174 265084
rect 196250 265072 196256 265084
rect 196308 265072 196314 265124
rect 170398 265004 170404 265056
rect 170456 265044 170462 265056
rect 170674 265044 170680 265056
rect 170456 265016 170680 265044
rect 170456 265004 170462 265016
rect 170674 265004 170680 265016
rect 170732 265044 170738 265056
rect 197906 265044 197912 265056
rect 170732 265016 197912 265044
rect 170732 265004 170738 265016
rect 197906 265004 197912 265016
rect 197964 265004 197970 265056
rect 119706 264936 119712 264988
rect 119764 264976 119770 264988
rect 152182 264976 152188 264988
rect 119764 264948 152188 264976
rect 119764 264936 119770 264948
rect 152182 264936 152188 264948
rect 152240 264976 152246 264988
rect 152458 264976 152464 264988
rect 152240 264948 152464 264976
rect 152240 264936 152246 264948
rect 152458 264936 152464 264948
rect 152516 264936 152522 264988
rect 160830 264936 160836 264988
rect 160888 264976 160894 264988
rect 193398 264976 193404 264988
rect 160888 264948 193404 264976
rect 160888 264936 160894 264948
rect 193398 264936 193404 264948
rect 193456 264936 193462 264988
rect 149698 264324 149704 264376
rect 149756 264364 149762 264376
rect 173434 264364 173440 264376
rect 149756 264336 173440 264364
rect 149756 264324 149762 264336
rect 173434 264324 173440 264336
rect 173492 264324 173498 264376
rect 139394 264256 139400 264308
rect 139452 264296 139458 264308
rect 178678 264296 178684 264308
rect 139452 264268 178684 264296
rect 139452 264256 139458 264268
rect 178678 264256 178684 264268
rect 178736 264256 178742 264308
rect 106918 264188 106924 264240
rect 106976 264228 106982 264240
rect 158714 264228 158720 264240
rect 106976 264200 158720 264228
rect 106976 264188 106982 264200
rect 158714 264188 158720 264200
rect 158772 264188 158778 264240
rect 119890 264052 119896 264104
rect 119948 264092 119954 264104
rect 137830 264092 137836 264104
rect 119948 264064 137836 264092
rect 119948 264052 119954 264064
rect 137830 264052 137836 264064
rect 137888 264052 137894 264104
rect 116762 263984 116768 264036
rect 116820 264024 116826 264036
rect 134426 264024 134432 264036
rect 116820 263996 134432 264024
rect 116820 263984 116826 263996
rect 134426 263984 134432 263996
rect 134484 264024 134490 264036
rect 134610 264024 134616 264036
rect 134484 263996 134616 264024
rect 134484 263984 134490 263996
rect 134610 263984 134616 263996
rect 134668 263984 134674 264036
rect 119522 263916 119528 263968
rect 119580 263956 119586 263968
rect 139394 263956 139400 263968
rect 119580 263928 139400 263956
rect 119580 263916 119586 263928
rect 139394 263916 139400 263928
rect 139452 263916 139458 263968
rect 112714 263848 112720 263900
rect 112772 263888 112778 263900
rect 133138 263888 133144 263900
rect 112772 263860 133144 263888
rect 112772 263848 112778 263860
rect 133138 263848 133144 263860
rect 133196 263848 133202 263900
rect 120902 263780 120908 263832
rect 120960 263820 120966 263832
rect 141418 263820 141424 263832
rect 120960 263792 141424 263820
rect 120960 263780 120966 263792
rect 141418 263780 141424 263792
rect 141476 263780 141482 263832
rect 119614 263712 119620 263764
rect 119672 263752 119678 263764
rect 142614 263752 142620 263764
rect 119672 263724 142620 263752
rect 119672 263712 119678 263724
rect 142614 263712 142620 263724
rect 142672 263712 142678 263764
rect 114002 263644 114008 263696
rect 114060 263684 114066 263696
rect 137186 263684 137192 263696
rect 114060 263656 137192 263684
rect 114060 263644 114066 263656
rect 137186 263644 137192 263656
rect 137244 263644 137250 263696
rect 173158 263644 173164 263696
rect 173216 263684 173222 263696
rect 173434 263684 173440 263696
rect 173216 263656 173440 263684
rect 173216 263644 173222 263656
rect 173434 263644 173440 263656
rect 173492 263684 173498 263696
rect 194962 263684 194968 263696
rect 173492 263656 194968 263684
rect 173492 263644 173498 263656
rect 194962 263644 194968 263656
rect 195020 263644 195026 263696
rect 120994 263576 121000 263628
rect 121052 263616 121058 263628
rect 151078 263616 151084 263628
rect 121052 263588 151084 263616
rect 121052 263576 121058 263588
rect 151078 263576 151084 263588
rect 151136 263576 151142 263628
rect 158714 263576 158720 263628
rect 158772 263616 158778 263628
rect 159358 263616 159364 263628
rect 158772 263588 159364 263616
rect 158772 263576 158778 263588
rect 159358 263576 159364 263588
rect 159416 263616 159422 263628
rect 190914 263616 190920 263628
rect 159416 263588 190920 263616
rect 159416 263576 159422 263588
rect 190914 263576 190920 263588
rect 190972 263576 190978 263628
rect 137462 263508 137468 263560
rect 137520 263548 137526 263560
rect 580258 263548 580264 263560
rect 137520 263520 580264 263548
rect 137520 263508 137526 263520
rect 580258 263508 580264 263520
rect 580316 263508 580322 263560
rect 147674 263440 147680 263492
rect 147732 263480 147738 263492
rect 148042 263480 148048 263492
rect 147732 263452 148048 263480
rect 147732 263440 147738 263452
rect 148042 263440 148048 263452
rect 148100 263440 148106 263492
rect 191006 263440 191012 263492
rect 191064 263480 191070 263492
rect 282914 263480 282920 263492
rect 191064 263452 282920 263480
rect 191064 263440 191070 263452
rect 282914 263440 282920 263452
rect 282972 263440 282978 263492
rect 191834 263372 191840 263424
rect 191892 263412 191898 263424
rect 218054 263412 218060 263424
rect 191892 263384 218060 263412
rect 191892 263372 191898 263384
rect 218054 263372 218060 263384
rect 218112 263372 218118 263424
rect 3510 263100 3516 263152
rect 3568 263140 3574 263152
rect 176746 263140 176752 263152
rect 3568 263112 176752 263140
rect 3568 263100 3574 263112
rect 176746 263100 176752 263112
rect 176804 263100 176810 263152
rect 179230 263100 179236 263152
rect 179288 263140 179294 263152
rect 192478 263140 192484 263152
rect 179288 263112 192484 263140
rect 179288 263100 179294 263112
rect 192478 263100 192484 263112
rect 192536 263100 192542 263152
rect 132034 263032 132040 263084
rect 132092 263072 132098 263084
rect 580350 263072 580356 263084
rect 132092 263044 580356 263072
rect 132092 263032 132098 263044
rect 580350 263032 580356 263044
rect 580408 263032 580414 263084
rect 167822 262964 167828 263016
rect 167880 263004 167886 263016
rect 192294 263004 192300 263016
rect 167880 262976 192300 263004
rect 167880 262964 167886 262976
rect 192294 262964 192300 262976
rect 192352 262964 192358 263016
rect 116670 262896 116676 262948
rect 116728 262936 116734 262948
rect 127618 262936 127624 262948
rect 116728 262908 127624 262936
rect 116728 262896 116734 262908
rect 127618 262896 127624 262908
rect 127676 262896 127682 262948
rect 131114 262896 131120 262948
rect 131172 262936 131178 262948
rect 131758 262936 131764 262948
rect 131172 262908 131764 262936
rect 131172 262896 131178 262908
rect 131758 262896 131764 262908
rect 131816 262936 131822 262948
rect 580442 262936 580448 262948
rect 131816 262908 580448 262936
rect 131816 262896 131822 262908
rect 580442 262896 580448 262908
rect 580500 262896 580506 262948
rect 3418 262828 3424 262880
rect 3476 262868 3482 262880
rect 178402 262868 178408 262880
rect 3476 262840 178408 262868
rect 3476 262828 3482 262840
rect 178402 262828 178408 262840
rect 178460 262828 178466 262880
rect 347774 262868 347780 262880
rect 195946 262840 347780 262868
rect 112530 262760 112536 262812
rect 112588 262800 112594 262812
rect 131114 262800 131120 262812
rect 112588 262772 131120 262800
rect 112588 262760 112594 262772
rect 131114 262760 131120 262772
rect 131172 262760 131178 262812
rect 166258 262760 166264 262812
rect 166316 262800 166322 262812
rect 192202 262800 192208 262812
rect 166316 262772 192208 262800
rect 166316 262760 166322 262772
rect 192202 262760 192208 262772
rect 192260 262760 192266 262812
rect 113726 262692 113732 262744
rect 113784 262732 113790 262744
rect 134518 262732 134524 262744
rect 113784 262704 134524 262732
rect 113784 262692 113790 262704
rect 134518 262692 134524 262704
rect 134576 262732 134582 262744
rect 134794 262732 134800 262744
rect 134576 262704 134800 262732
rect 134576 262692 134582 262704
rect 134794 262692 134800 262704
rect 134852 262692 134858 262744
rect 153194 262692 153200 262744
rect 153252 262732 153258 262744
rect 158714 262732 158720 262744
rect 153252 262704 158720 262732
rect 153252 262692 153258 262704
rect 158714 262692 158720 262704
rect 158772 262692 158778 262744
rect 164970 262692 164976 262744
rect 165028 262732 165034 262744
rect 193582 262732 193588 262744
rect 165028 262704 193588 262732
rect 165028 262692 165034 262704
rect 193582 262692 193588 262704
rect 193640 262692 193646 262744
rect 116578 262624 116584 262676
rect 116636 262664 116642 262676
rect 131114 262664 131120 262676
rect 116636 262636 131120 262664
rect 116636 262624 116642 262636
rect 131114 262624 131120 262636
rect 131172 262624 131178 262676
rect 153838 262624 153844 262676
rect 153896 262664 153902 262676
rect 188246 262664 188252 262676
rect 153896 262636 188252 262664
rect 153896 262624 153902 262636
rect 188246 262624 188252 262636
rect 188304 262664 188310 262676
rect 195946 262664 195974 262840
rect 347774 262828 347780 262840
rect 347832 262828 347838 262880
rect 188304 262636 195974 262664
rect 188304 262624 188310 262636
rect 116486 262556 116492 262608
rect 116544 262596 116550 262608
rect 144178 262596 144184 262608
rect 116544 262568 144184 262596
rect 116544 262556 116550 262568
rect 144178 262556 144184 262568
rect 144236 262556 144242 262608
rect 155862 262556 155868 262608
rect 155920 262596 155926 262608
rect 191006 262596 191012 262608
rect 155920 262568 191012 262596
rect 155920 262556 155926 262568
rect 191006 262556 191012 262568
rect 191064 262556 191070 262608
rect 113910 262488 113916 262540
rect 113968 262528 113974 262540
rect 142246 262528 142252 262540
rect 113968 262500 142252 262528
rect 113968 262488 113974 262500
rect 142246 262488 142252 262500
rect 142304 262528 142310 262540
rect 142890 262528 142896 262540
rect 142304 262500 142896 262528
rect 142304 262488 142310 262500
rect 142890 262488 142896 262500
rect 142948 262488 142954 262540
rect 157150 262488 157156 262540
rect 157208 262528 157214 262540
rect 191834 262528 191840 262540
rect 157208 262500 191840 262528
rect 157208 262488 157214 262500
rect 191834 262488 191840 262500
rect 191892 262488 191898 262540
rect 118418 262420 118424 262472
rect 118476 262460 118482 262472
rect 125962 262460 125968 262472
rect 118476 262432 125968 262460
rect 118476 262420 118482 262432
rect 125962 262420 125968 262432
rect 126020 262420 126026 262472
rect 181806 262420 181812 262472
rect 181864 262460 181870 262472
rect 196342 262460 196348 262472
rect 181864 262432 196348 262460
rect 181864 262420 181870 262432
rect 196342 262420 196348 262432
rect 196400 262420 196406 262472
rect 118234 262352 118240 262404
rect 118292 262392 118298 262404
rect 129274 262392 129280 262404
rect 118292 262364 129280 262392
rect 118292 262352 118298 262364
rect 129274 262352 129280 262364
rect 129332 262352 129338 262404
rect 182910 262352 182916 262404
rect 182968 262392 182974 262404
rect 190546 262392 190552 262404
rect 182968 262364 190552 262392
rect 182968 262352 182974 262364
rect 190546 262352 190552 262364
rect 190604 262352 190610 262404
rect 181254 262284 181260 262336
rect 181312 262324 181318 262336
rect 190638 262324 190644 262336
rect 181312 262296 190644 262324
rect 181312 262284 181318 262296
rect 190638 262284 190644 262296
rect 190696 262284 190702 262336
rect 116854 262216 116860 262268
rect 116912 262256 116918 262268
rect 122742 262256 122748 262268
rect 116912 262228 122748 262256
rect 116912 262216 116918 262228
rect 122742 262216 122748 262228
rect 122800 262216 122806 262268
rect 184566 262216 184572 262268
rect 184624 262256 184630 262268
rect 189166 262256 189172 262268
rect 184624 262228 189172 262256
rect 184624 262216 184630 262228
rect 189166 262216 189172 262228
rect 189224 262216 189230 262268
rect 129826 261536 129832 261588
rect 129884 261576 129890 261588
rect 189718 261576 189724 261588
rect 129884 261548 189724 261576
rect 129884 261536 129890 261548
rect 189718 261536 189724 261548
rect 189776 261536 189782 261588
rect 178402 261468 178408 261520
rect 178460 261508 178466 261520
rect 200574 261508 200580 261520
rect 178460 261480 200580 261508
rect 178460 261468 178466 261480
rect 200574 261468 200580 261480
rect 200632 261468 200638 261520
rect 131114 261400 131120 261452
rect 131172 261440 131178 261452
rect 471238 261440 471244 261452
rect 131172 261412 471244 261440
rect 131172 261400 131178 261412
rect 471238 261400 471244 261412
rect 471296 261400 471302 261452
rect 118326 261332 118332 261384
rect 118384 261372 118390 261384
rect 127342 261372 127348 261384
rect 118384 261344 127348 261372
rect 118384 261332 118390 261344
rect 127342 261332 127348 261344
rect 127400 261332 127406 261384
rect 183462 261332 183468 261384
rect 183520 261372 183526 261384
rect 197814 261372 197820 261384
rect 183520 261344 197820 261372
rect 183520 261332 183526 261344
rect 197814 261332 197820 261344
rect 197872 261332 197878 261384
rect 14458 261264 14464 261316
rect 14516 261304 14522 261316
rect 176194 261304 176200 261316
rect 14516 261276 176200 261304
rect 14516 261264 14522 261276
rect 176194 261264 176200 261276
rect 176252 261264 176258 261316
rect 177298 261264 177304 261316
rect 177356 261304 177362 261316
rect 193766 261304 193772 261316
rect 177356 261276 193772 261304
rect 177356 261264 177362 261276
rect 193766 261264 193772 261276
rect 193824 261264 193830 261316
rect 111242 261196 111248 261248
rect 111300 261236 111306 261248
rect 134334 261236 134340 261248
rect 111300 261208 134340 261236
rect 111300 261196 111306 261208
rect 134334 261196 134340 261208
rect 134392 261196 134398 261248
rect 180518 261196 180524 261248
rect 180576 261236 180582 261248
rect 199286 261236 199292 261248
rect 180576 261208 199292 261236
rect 180576 261196 180582 261208
rect 199286 261196 199292 261208
rect 199344 261196 199350 261248
rect 117958 261128 117964 261180
rect 118016 261168 118022 261180
rect 127066 261168 127072 261180
rect 118016 261140 127072 261168
rect 118016 261128 118022 261140
rect 127066 261128 127072 261140
rect 127124 261128 127130 261180
rect 127342 261128 127348 261180
rect 127400 261168 127406 261180
rect 132862 261168 132868 261180
rect 127400 261140 132868 261168
rect 127400 261128 127406 261140
rect 132862 261128 132868 261140
rect 132920 261128 132926 261180
rect 176746 261128 176752 261180
rect 176804 261168 176810 261180
rect 196710 261168 196716 261180
rect 176804 261140 196716 261168
rect 176804 261128 176810 261140
rect 196710 261128 196716 261140
rect 196768 261128 196774 261180
rect 110874 261060 110880 261112
rect 110932 261100 110938 261112
rect 128722 261100 128728 261112
rect 110932 261072 128728 261100
rect 110932 261060 110938 261072
rect 128722 261060 128728 261072
rect 128780 261060 128786 261112
rect 158714 261060 158720 261112
rect 158772 261100 158778 261112
rect 193674 261100 193680 261112
rect 158772 261072 193680 261100
rect 158772 261060 158778 261072
rect 193674 261060 193680 261072
rect 193732 261060 193738 261112
rect 111058 260992 111064 261044
rect 111116 261032 111122 261044
rect 130378 261032 130384 261044
rect 111116 261004 130384 261032
rect 111116 260992 111122 261004
rect 130378 260992 130384 261004
rect 130436 260992 130442 261044
rect 181990 260992 181996 261044
rect 182048 261032 182054 261044
rect 200482 261032 200488 261044
rect 182048 261004 200488 261032
rect 182048 260992 182054 261004
rect 200482 260992 200488 261004
rect 200540 260992 200546 261044
rect 176194 260924 176200 260976
rect 176252 260964 176258 260976
rect 195054 260964 195060 260976
rect 176252 260936 195060 260964
rect 176252 260924 176258 260936
rect 195054 260924 195060 260936
rect 195112 260924 195118 260976
rect 114094 260856 114100 260908
rect 114152 260896 114158 260908
rect 125594 260896 125600 260908
rect 114152 260868 125600 260896
rect 114152 260856 114158 260868
rect 125594 260856 125600 260868
rect 125652 260856 125658 260908
rect 184014 260856 184020 260908
rect 184072 260896 184078 260908
rect 199194 260896 199200 260908
rect 184072 260868 199200 260896
rect 184072 260856 184078 260868
rect 199194 260856 199200 260868
rect 199252 260856 199258 260908
rect 120810 260788 120816 260840
rect 120868 260828 120874 260840
rect 123202 260828 123208 260840
rect 120868 260800 123208 260828
rect 120868 260788 120874 260800
rect 123202 260788 123208 260800
rect 123260 260788 123266 260840
rect 119798 260720 119804 260772
rect 119856 260760 119862 260772
rect 122834 260760 122840 260772
rect 119856 260732 122840 260760
rect 119856 260720 119862 260732
rect 122834 260720 122840 260732
rect 122892 260720 122898 260772
rect 122742 260652 122748 260704
rect 122800 260692 122806 260704
rect 124306 260692 124312 260704
rect 122800 260664 124312 260692
rect 122800 260652 122806 260664
rect 124306 260652 124312 260664
rect 124364 260652 124370 260704
rect 173894 260448 173900 260500
rect 173952 260488 173958 260500
rect 193490 260488 193496 260500
rect 173952 260460 193496 260488
rect 173952 260448 173958 260460
rect 193490 260448 193496 260460
rect 193548 260448 193554 260500
rect 134334 260380 134340 260432
rect 134392 260420 134398 260432
rect 188982 260420 188988 260432
rect 134392 260392 188988 260420
rect 134392 260380 134398 260392
rect 188982 260380 188988 260392
rect 189040 260380 189046 260432
rect 4798 260312 4804 260364
rect 4856 260352 4862 260364
rect 177298 260352 177304 260364
rect 4856 260324 177304 260352
rect 4856 260312 4862 260324
rect 177298 260312 177304 260324
rect 177356 260312 177362 260364
rect 175918 260244 175924 260296
rect 175976 260284 175982 260296
rect 192386 260284 192392 260296
rect 175976 260256 192392 260284
rect 175976 260244 175982 260256
rect 192386 260244 192392 260256
rect 192444 260244 192450 260296
rect 135254 260176 135260 260228
rect 135312 260216 135318 260228
rect 136220 260216 136226 260228
rect 135312 260188 136226 260216
rect 135312 260176 135318 260188
rect 136220 260176 136226 260188
rect 136278 260176 136284 260228
rect 155954 260176 155960 260228
rect 156012 260216 156018 260228
rect 156644 260216 156650 260228
rect 156012 260188 156650 260216
rect 156012 260176 156018 260188
rect 156644 260176 156650 260188
rect 156702 260176 156708 260228
rect 166994 260176 167000 260228
rect 167052 260216 167058 260228
rect 167684 260216 167690 260228
rect 167052 260188 167690 260216
rect 167052 260176 167058 260188
rect 167684 260176 167690 260188
rect 167742 260176 167748 260228
rect 169754 260176 169760 260228
rect 169812 260216 169818 260228
rect 170996 260216 171002 260228
rect 169812 260188 171002 260216
rect 169812 260176 169818 260188
rect 170996 260176 171002 260188
rect 171054 260176 171060 260228
rect 191190 260216 191196 260228
rect 171106 260188 191196 260216
rect 169202 260108 169208 260160
rect 169260 260148 169266 260160
rect 171106 260148 171134 260188
rect 191190 260176 191196 260188
rect 191248 260176 191254 260228
rect 169260 260120 171134 260148
rect 169260 260108 169266 260120
rect 167684 260040 167690 260092
rect 167742 260080 167748 260092
rect 189626 260080 189632 260092
rect 167742 260052 189632 260080
rect 167742 260040 167748 260052
rect 189626 260040 189632 260052
rect 189684 260040 189690 260092
rect 112622 259972 112628 260024
rect 112680 260012 112686 260024
rect 123754 260012 123760 260024
rect 112680 259984 123760 260012
rect 112680 259972 112686 259984
rect 123754 259972 123760 259984
rect 123812 259972 123818 260024
rect 164694 259972 164700 260024
rect 164752 260012 164758 260024
rect 189534 260012 189540 260024
rect 164752 259984 189540 260012
rect 164752 259972 164758 259984
rect 189534 259972 189540 259984
rect 189592 259972 189598 260024
rect 118142 259904 118148 259956
rect 118200 259944 118206 259956
rect 135254 259944 135260 259956
rect 118200 259916 135260 259944
rect 118200 259904 118206 259916
rect 135254 259904 135260 259916
rect 135312 259904 135318 259956
rect 166166 259904 166172 259956
rect 166224 259944 166230 259956
rect 191006 259944 191012 259956
rect 166224 259916 191012 259944
rect 166224 259904 166230 259916
rect 191006 259904 191012 259916
rect 191064 259904 191070 259956
rect 119338 259836 119344 259888
rect 119396 259876 119402 259888
rect 149146 259876 149152 259888
rect 119396 259848 149152 259876
rect 119396 259836 119402 259848
rect 149146 259836 149152 259848
rect 149204 259836 149210 259888
rect 156966 259836 156972 259888
rect 157024 259876 157030 259888
rect 189350 259876 189356 259888
rect 157024 259848 189356 259876
rect 157024 259836 157030 259848
rect 189350 259836 189356 259848
rect 189408 259836 189414 259888
rect 118050 259768 118056 259820
rect 118108 259808 118114 259820
rect 150434 259808 150440 259820
rect 118108 259780 150440 259808
rect 118108 259768 118114 259780
rect 150434 259768 150440 259780
rect 150492 259808 150498 259820
rect 151354 259808 151360 259820
rect 150492 259780 151360 259808
rect 150492 259768 150498 259780
rect 151354 259768 151360 259780
rect 151412 259768 151418 259820
rect 171134 259768 171140 259820
rect 171192 259808 171198 259820
rect 203242 259808 203248 259820
rect 171192 259780 203248 259808
rect 171192 259768 171198 259780
rect 203242 259768 203248 259780
rect 203300 259768 203306 259820
rect 119430 259700 119436 259752
rect 119488 259740 119494 259752
rect 153194 259740 153200 259752
rect 119488 259712 153200 259740
rect 119488 259700 119494 259712
rect 153194 259700 153200 259712
rect 153252 259700 153258 259752
rect 158070 259700 158076 259752
rect 158128 259740 158134 259752
rect 191098 259740 191104 259752
rect 158128 259712 191104 259740
rect 158128 259700 158134 259712
rect 191098 259700 191104 259712
rect 191156 259700 191162 259752
rect 115290 259632 115296 259684
rect 115348 259672 115354 259684
rect 128354 259672 128360 259684
rect 115348 259644 128360 259672
rect 115348 259632 115354 259644
rect 128354 259632 128360 259644
rect 128412 259632 128418 259684
rect 184934 259632 184940 259684
rect 184992 259672 184998 259684
rect 196618 259672 196624 259684
rect 184992 259644 196624 259672
rect 184992 259632 184998 259644
rect 196618 259632 196624 259644
rect 196676 259632 196682 259684
rect 117866 259564 117872 259616
rect 117924 259604 117930 259616
rect 178034 259604 178040 259616
rect 117924 259576 178040 259604
rect 117924 259564 117930 259576
rect 178034 259564 178040 259576
rect 178092 259604 178098 259616
rect 195238 259604 195244 259616
rect 178092 259576 195244 259604
rect 178092 259564 178098 259576
rect 195238 259564 195244 259576
rect 195296 259564 195302 259616
rect 115474 259496 115480 259548
rect 115532 259536 115538 259548
rect 126514 259536 126520 259548
rect 115532 259508 126520 259536
rect 115532 259496 115538 259508
rect 126514 259496 126520 259508
rect 126572 259496 126578 259548
rect 180150 259496 180156 259548
rect 180208 259536 180214 259548
rect 197722 259536 197728 259548
rect 180208 259508 197728 259536
rect 180208 259496 180214 259508
rect 197722 259496 197728 259508
rect 197780 259496 197786 259548
rect 120718 259428 120724 259480
rect 120776 259468 120782 259480
rect 124858 259468 124864 259480
rect 120776 259440 124864 259468
rect 120776 259428 120782 259440
rect 124858 259428 124864 259440
rect 124916 259428 124922 259480
rect 133230 259428 133236 259480
rect 133288 259468 133294 259480
rect 472618 259468 472624 259480
rect 133288 259440 472624 259468
rect 133288 259428 133294 259440
rect 472618 259428 472624 259440
rect 472676 259428 472682 259480
rect 188982 259360 188988 259412
rect 189040 259400 189046 259412
rect 580166 259400 580172 259412
rect 189040 259372 580172 259400
rect 189040 259360 189046 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 472618 245556 472624 245608
rect 472676 245596 472682 245608
rect 580166 245596 580172 245608
rect 472676 245568 580172 245596
rect 472676 245556 472682 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 14458 241448 14464 241460
rect 3568 241420 14464 241448
rect 3568 241408 3574 241420
rect 14458 241408 14464 241420
rect 14516 241408 14522 241460
rect 2774 215228 2780 215280
rect 2832 215268 2838 215280
rect 4798 215268 4804 215280
rect 2832 215240 4804 215268
rect 2832 215228 2838 215240
rect 4798 215228 4804 215240
rect 4856 215228 4862 215280
rect 471238 206932 471244 206984
rect 471296 206972 471302 206984
rect 579798 206972 579804 206984
rect 471296 206944 579804 206972
rect 471296 206932 471302 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 190454 200784 190460 200796
rect 128924 200756 131712 200784
rect 128924 200728 128952 200756
rect 131684 200728 131712 200756
rect 178788 200756 190460 200784
rect 178788 200728 178816 200756
rect 190454 200744 190460 200756
rect 190512 200744 190518 200796
rect 128906 200676 128912 200728
rect 128964 200676 128970 200728
rect 129274 200676 129280 200728
rect 129332 200716 129338 200728
rect 131574 200716 131580 200728
rect 129332 200688 131580 200716
rect 129332 200676 129338 200688
rect 131574 200676 131580 200688
rect 131632 200676 131638 200728
rect 131666 200676 131672 200728
rect 131724 200676 131730 200728
rect 178770 200676 178776 200728
rect 178828 200676 178834 200728
rect 132218 200648 132224 200660
rect 125566 200620 132224 200648
rect 111610 200540 111616 200592
rect 111668 200580 111674 200592
rect 125566 200580 125594 200620
rect 132218 200608 132224 200620
rect 132276 200608 132282 200660
rect 172486 200620 173894 200648
rect 111668 200552 125594 200580
rect 111668 200540 111674 200552
rect 128078 200540 128084 200592
rect 128136 200580 128142 200592
rect 131942 200580 131948 200592
rect 128136 200552 131948 200580
rect 128136 200540 128142 200552
rect 131942 200540 131948 200552
rect 132000 200540 132006 200592
rect 132034 200540 132040 200592
rect 132092 200580 132098 200592
rect 172486 200580 172514 200620
rect 132092 200552 138014 200580
rect 132092 200540 132098 200552
rect 108942 200472 108948 200524
rect 109000 200512 109006 200524
rect 131758 200512 131764 200524
rect 109000 200484 131764 200512
rect 109000 200472 109006 200484
rect 131758 200472 131764 200484
rect 131816 200472 131822 200524
rect 137986 200512 138014 200552
rect 159422 200552 172514 200580
rect 173866 200580 173894 200620
rect 173866 200552 179414 200580
rect 137986 200484 151170 200512
rect 130470 200404 130476 200456
rect 130528 200444 130534 200456
rect 131850 200444 131856 200456
rect 130528 200416 131856 200444
rect 130528 200404 130534 200416
rect 131850 200404 131856 200416
rect 131908 200404 131914 200456
rect 137986 200416 149606 200444
rect 123938 200336 123944 200388
rect 123996 200376 124002 200388
rect 137986 200376 138014 200416
rect 123996 200348 138014 200376
rect 139366 200348 148502 200376
rect 123996 200336 124002 200348
rect 121086 200268 121092 200320
rect 121144 200308 121150 200320
rect 139366 200308 139394 200348
rect 121144 200280 139394 200308
rect 121144 200268 121150 200280
rect 131482 200200 131488 200252
rect 131540 200240 131546 200252
rect 131540 200212 147398 200240
rect 131540 200200 131546 200212
rect 131758 200132 131764 200184
rect 131816 200172 131822 200184
rect 131816 200144 137002 200172
rect 131816 200132 131822 200144
rect 131850 200064 131856 200116
rect 131908 200104 131914 200116
rect 131908 200076 136910 200104
rect 131908 200064 131914 200076
rect 129090 199928 129096 199980
rect 129148 199968 129154 199980
rect 132218 199968 132224 199980
rect 129148 199940 132224 199968
rect 129148 199928 129154 199940
rect 132218 199928 132224 199940
rect 132276 199928 132282 199980
rect 132328 199940 132678 199968
rect 128354 199860 128360 199912
rect 128412 199900 128418 199912
rect 132328 199900 132356 199940
rect 132650 199912 132678 199940
rect 132834 199940 134058 199968
rect 132540 199900 132546 199912
rect 128412 199872 132356 199900
rect 132466 199872 132546 199900
rect 128412 199860 128418 199872
rect 128538 199792 128544 199844
rect 128596 199832 128602 199844
rect 132126 199832 132132 199844
rect 128596 199804 132132 199832
rect 128596 199792 128602 199804
rect 132126 199792 132132 199804
rect 132184 199792 132190 199844
rect 131758 199724 131764 199776
rect 131816 199764 131822 199776
rect 132466 199764 132494 199872
rect 132540 199860 132546 199872
rect 132598 199860 132604 199912
rect 132632 199860 132638 199912
rect 132690 199860 132696 199912
rect 131816 199736 132494 199764
rect 131816 199724 131822 199736
rect 126146 199656 126152 199708
rect 126204 199696 126210 199708
rect 132834 199696 132862 199940
rect 134030 199912 134058 199940
rect 134490 199940 134886 199968
rect 133000 199860 133006 199912
rect 133058 199860 133064 199912
rect 133184 199860 133190 199912
rect 133242 199860 133248 199912
rect 133736 199860 133742 199912
rect 133794 199860 133800 199912
rect 134012 199860 134018 199912
rect 134070 199860 134076 199912
rect 134380 199860 134386 199912
rect 134438 199860 134444 199912
rect 133018 199832 133046 199860
rect 126204 199668 132862 199696
rect 132926 199804 133046 199832
rect 126204 199656 126210 199668
rect 118510 199588 118516 199640
rect 118568 199628 118574 199640
rect 131850 199628 131856 199640
rect 118568 199600 131856 199628
rect 118568 199588 118574 199600
rect 131850 199588 131856 199600
rect 131908 199588 131914 199640
rect 131942 199588 131948 199640
rect 132000 199628 132006 199640
rect 132926 199628 132954 199804
rect 133202 199640 133230 199860
rect 133754 199776 133782 199860
rect 133690 199724 133696 199776
rect 133748 199736 133782 199776
rect 133748 199724 133754 199736
rect 133966 199724 133972 199776
rect 134024 199764 134030 199776
rect 134398 199764 134426 199860
rect 134024 199736 134426 199764
rect 134024 199724 134030 199736
rect 134490 199640 134518 199940
rect 134564 199860 134570 199912
rect 134622 199860 134628 199912
rect 134582 199696 134610 199860
rect 134858 199844 134886 199940
rect 136330 199940 136818 199968
rect 136330 199912 136358 199940
rect 135024 199860 135030 199912
rect 135082 199860 135088 199912
rect 135392 199860 135398 199912
rect 135450 199860 135456 199912
rect 135576 199860 135582 199912
rect 135634 199860 135640 199912
rect 135668 199860 135674 199912
rect 135726 199860 135732 199912
rect 135760 199860 135766 199912
rect 135818 199900 135824 199912
rect 135818 199872 135944 199900
rect 135818 199860 135824 199872
rect 134840 199792 134846 199844
rect 134898 199792 134904 199844
rect 134582 199668 134702 199696
rect 132000 199600 132954 199628
rect 132000 199588 132006 199600
rect 133138 199588 133144 199640
rect 133196 199600 133230 199640
rect 133196 199588 133202 199600
rect 134426 199588 134432 199640
rect 134484 199600 134518 199640
rect 134484 199588 134490 199600
rect 117038 199520 117044 199572
rect 117096 199560 117102 199572
rect 131482 199560 131488 199572
rect 117096 199532 131488 199560
rect 117096 199520 117102 199532
rect 131482 199520 131488 199532
rect 131540 199520 131546 199572
rect 115658 199452 115664 199504
rect 115716 199492 115722 199504
rect 132954 199492 132960 199504
rect 115716 199464 132960 199492
rect 115716 199452 115722 199464
rect 132954 199452 132960 199464
rect 133012 199452 133018 199504
rect 133874 199452 133880 199504
rect 133932 199492 133938 199504
rect 134334 199492 134340 199504
rect 133932 199464 134340 199492
rect 133932 199452 133938 199464
rect 134334 199452 134340 199464
rect 134392 199452 134398 199504
rect 115750 199384 115756 199436
rect 115808 199424 115814 199436
rect 132494 199424 132500 199436
rect 115808 199396 132500 199424
rect 115808 199384 115814 199396
rect 132494 199384 132500 199396
rect 132552 199384 132558 199436
rect 134674 199368 134702 199668
rect 135042 199640 135070 199860
rect 135300 199792 135306 199844
rect 135358 199792 135364 199844
rect 134978 199588 134984 199640
rect 135036 199600 135070 199640
rect 135036 199588 135042 199600
rect 134794 199452 134800 199504
rect 134852 199492 134858 199504
rect 135318 199492 135346 199792
rect 135410 199560 135438 199860
rect 135594 199708 135622 199860
rect 135686 199776 135714 199860
rect 135686 199736 135720 199776
rect 135714 199724 135720 199736
rect 135772 199724 135778 199776
rect 135594 199668 135628 199708
rect 135622 199656 135628 199668
rect 135680 199656 135686 199708
rect 135916 199640 135944 199872
rect 136036 199860 136042 199912
rect 136094 199900 136100 199912
rect 136094 199860 136128 199900
rect 136220 199860 136226 199912
rect 136278 199860 136284 199912
rect 136312 199860 136318 199912
rect 136370 199860 136376 199912
rect 135898 199588 135904 199640
rect 135956 199588 135962 199640
rect 136100 199628 136128 199860
rect 136238 199776 136266 199860
rect 136790 199832 136818 199940
rect 136882 199912 136910 200076
rect 136974 200036 137002 200144
rect 136974 200008 138842 200036
rect 138814 199912 138842 200008
rect 138998 200008 142246 200036
rect 136864 199860 136870 199912
rect 136922 199860 136928 199912
rect 136956 199860 136962 199912
rect 137014 199860 137020 199912
rect 137140 199900 137146 199912
rect 137066 199872 137146 199900
rect 136790 199804 136864 199832
rect 136238 199736 136272 199776
rect 136266 199724 136272 199736
rect 136324 199724 136330 199776
rect 136634 199628 136640 199640
rect 136100 199600 136640 199628
rect 136634 199588 136640 199600
rect 136692 199588 136698 199640
rect 135530 199560 135536 199572
rect 135410 199532 135536 199560
rect 135530 199520 135536 199532
rect 135588 199520 135594 199572
rect 136542 199520 136548 199572
rect 136600 199560 136606 199572
rect 136836 199560 136864 199804
rect 136974 199776 137002 199860
rect 136910 199724 136916 199776
rect 136968 199736 137002 199776
rect 136968 199724 136974 199736
rect 137066 199708 137094 199872
rect 137140 199860 137146 199872
rect 137198 199860 137204 199912
rect 137416 199900 137422 199912
rect 137388 199860 137422 199900
rect 137474 199860 137480 199912
rect 137508 199860 137514 199912
rect 137566 199860 137572 199912
rect 137600 199860 137606 199912
rect 137658 199860 137664 199912
rect 138336 199860 138342 199912
rect 138394 199860 138400 199912
rect 138612 199860 138618 199912
rect 138670 199860 138676 199912
rect 138704 199860 138710 199912
rect 138762 199860 138768 199912
rect 138796 199860 138802 199912
rect 138854 199860 138860 199912
rect 138888 199860 138894 199912
rect 138946 199860 138952 199912
rect 137232 199832 137238 199844
rect 137204 199792 137238 199832
rect 137290 199792 137296 199844
rect 137204 199708 137232 199792
rect 137066 199668 137100 199708
rect 137094 199656 137100 199668
rect 137152 199656 137158 199708
rect 137186 199656 137192 199708
rect 137244 199656 137250 199708
rect 136600 199532 136864 199560
rect 136600 199520 136606 199532
rect 137278 199520 137284 199572
rect 137336 199560 137342 199572
rect 137388 199560 137416 199860
rect 137526 199776 137554 199860
rect 137462 199724 137468 199776
rect 137520 199736 137554 199776
rect 137520 199724 137526 199736
rect 137618 199640 137646 199860
rect 138354 199640 138382 199860
rect 138630 199708 138658 199860
rect 138722 199832 138750 199860
rect 138722 199804 138796 199832
rect 138768 199708 138796 199804
rect 138906 199776 138934 199860
rect 138842 199724 138848 199776
rect 138900 199736 138934 199776
rect 138900 199724 138906 199736
rect 138630 199668 138664 199708
rect 138658 199656 138664 199668
rect 138716 199656 138722 199708
rect 138750 199656 138756 199708
rect 138808 199656 138814 199708
rect 138998 199696 139026 200008
rect 139228 199940 141878 199968
rect 139072 199792 139078 199844
rect 139130 199832 139136 199844
rect 139130 199792 139164 199832
rect 138952 199668 139026 199696
rect 137618 199600 137652 199640
rect 137646 199588 137652 199600
rect 137704 199588 137710 199640
rect 138354 199600 138388 199640
rect 138382 199588 138388 199600
rect 138440 199588 138446 199640
rect 137336 199532 137416 199560
rect 137336 199520 137342 199532
rect 137922 199520 137928 199572
rect 137980 199560 137986 199572
rect 138952 199560 138980 199668
rect 137980 199532 138980 199560
rect 137980 199520 137986 199532
rect 139026 199520 139032 199572
rect 139084 199560 139090 199572
rect 139136 199560 139164 199792
rect 139228 199572 139256 199940
rect 141850 199912 141878 199940
rect 142218 199912 142246 200008
rect 142310 199940 143166 199968
rect 139716 199900 139722 199912
rect 139320 199872 139722 199900
rect 139084 199532 139164 199560
rect 139084 199520 139090 199532
rect 139210 199520 139216 199572
rect 139268 199520 139274 199572
rect 134852 199464 135346 199492
rect 134852 199452 134858 199464
rect 137554 199452 137560 199504
rect 137612 199492 137618 199504
rect 139320 199492 139348 199872
rect 139716 199860 139722 199872
rect 139774 199860 139780 199912
rect 139808 199860 139814 199912
rect 139866 199860 139872 199912
rect 139900 199860 139906 199912
rect 139958 199860 139964 199912
rect 139992 199860 139998 199912
rect 140050 199860 140056 199912
rect 140268 199860 140274 199912
rect 140326 199860 140332 199912
rect 140452 199860 140458 199912
rect 140510 199860 140516 199912
rect 140728 199860 140734 199912
rect 140786 199860 140792 199912
rect 141188 199860 141194 199912
rect 141246 199860 141252 199912
rect 141464 199860 141470 199912
rect 141522 199900 141528 199912
rect 141522 199872 141786 199900
rect 141522 199860 141528 199872
rect 139826 199708 139854 199860
rect 139762 199656 139768 199708
rect 139820 199668 139854 199708
rect 139820 199656 139826 199668
rect 139918 199640 139946 199860
rect 140010 199776 140038 199860
rect 140010 199736 140044 199776
rect 140038 199724 140044 199736
rect 140096 199724 140102 199776
rect 140286 199708 140314 199860
rect 140268 199656 140274 199708
rect 140326 199656 140332 199708
rect 139918 199600 139952 199640
rect 139946 199588 139952 199600
rect 140004 199588 140010 199640
rect 140470 199628 140498 199860
rect 140746 199640 140774 199860
rect 140590 199628 140596 199640
rect 140470 199600 140596 199628
rect 140590 199588 140596 199600
rect 140648 199588 140654 199640
rect 140746 199600 140780 199640
rect 140774 199588 140780 199600
rect 140832 199588 140838 199640
rect 141206 199628 141234 199860
rect 141648 199792 141654 199844
rect 141706 199792 141712 199844
rect 141666 199708 141694 199792
rect 141602 199656 141608 199708
rect 141660 199668 141694 199708
rect 141660 199656 141666 199668
rect 141418 199628 141424 199640
rect 141206 199600 141424 199628
rect 141418 199588 141424 199600
rect 141476 199588 141482 199640
rect 141758 199628 141786 199872
rect 141832 199860 141838 199912
rect 141890 199860 141896 199912
rect 141924 199860 141930 199912
rect 141982 199860 141988 199912
rect 142200 199860 142206 199912
rect 142258 199860 142264 199912
rect 141942 199776 141970 199860
rect 141878 199724 141884 199776
rect 141936 199736 141970 199776
rect 141936 199724 141942 199736
rect 142154 199724 142160 199776
rect 142212 199764 142218 199776
rect 142310 199764 142338 199940
rect 143138 199912 143166 199940
rect 144150 199940 144362 199968
rect 144150 199912 144178 199940
rect 142384 199860 142390 199912
rect 142442 199860 142448 199912
rect 142752 199900 142758 199912
rect 142586 199872 142758 199900
rect 142212 199736 142338 199764
rect 142212 199724 142218 199736
rect 142402 199640 142430 199860
rect 142062 199628 142068 199640
rect 141758 199600 142068 199628
rect 142062 199588 142068 199600
rect 142120 199588 142126 199640
rect 142402 199600 142436 199640
rect 142430 199588 142436 199600
rect 142488 199588 142494 199640
rect 137612 199464 139348 199492
rect 137612 199452 137618 199464
rect 140774 199452 140780 199504
rect 140832 199492 140838 199504
rect 141142 199492 141148 199504
rect 140832 199464 141148 199492
rect 140832 199452 140838 199464
rect 141142 199452 141148 199464
rect 141200 199452 141206 199504
rect 142586 199492 142614 199872
rect 142752 199860 142758 199872
rect 142810 199860 142816 199912
rect 143028 199860 143034 199912
rect 143086 199860 143092 199912
rect 143120 199860 143126 199912
rect 143178 199860 143184 199912
rect 143304 199860 143310 199912
rect 143362 199860 143368 199912
rect 143672 199860 143678 199912
rect 143730 199860 143736 199912
rect 143856 199860 143862 199912
rect 143914 199860 143920 199912
rect 143948 199860 143954 199912
rect 144006 199860 144012 199912
rect 144132 199860 144138 199912
rect 144190 199860 144196 199912
rect 144224 199860 144230 199912
rect 144282 199860 144288 199912
rect 142660 199792 142666 199844
rect 142718 199792 142724 199844
rect 142678 199708 142706 199792
rect 143046 199764 143074 199860
rect 143212 199792 143218 199844
rect 143270 199792 143276 199844
rect 143000 199736 143074 199764
rect 142678 199668 142712 199708
rect 142706 199656 142712 199668
rect 142764 199656 142770 199708
rect 143000 199572 143028 199736
rect 143074 199656 143080 199708
rect 143132 199696 143138 199708
rect 143230 199696 143258 199792
rect 143132 199668 143258 199696
rect 143132 199656 143138 199668
rect 143322 199640 143350 199860
rect 143690 199640 143718 199860
rect 143874 199832 143902 199860
rect 143828 199804 143902 199832
rect 143828 199640 143856 199804
rect 143966 199776 143994 199860
rect 143902 199724 143908 199776
rect 143960 199736 143994 199776
rect 143960 199724 143966 199736
rect 144242 199696 144270 199860
rect 144104 199668 144270 199696
rect 144104 199640 144132 199668
rect 143258 199588 143264 199640
rect 143316 199600 143350 199640
rect 143316 199588 143322 199600
rect 143626 199588 143632 199640
rect 143684 199600 143718 199640
rect 143684 199588 143690 199600
rect 143810 199588 143816 199640
rect 143868 199588 143874 199640
rect 144086 199588 144092 199640
rect 144144 199588 144150 199640
rect 144178 199588 144184 199640
rect 144236 199628 144242 199640
rect 144334 199628 144362 199940
rect 144564 199940 145006 199968
rect 144564 199640 144592 199940
rect 144978 199912 145006 199940
rect 145990 199940 146248 199968
rect 145990 199912 146018 199940
rect 144684 199860 144690 199912
rect 144742 199860 144748 199912
rect 144960 199860 144966 199912
rect 145018 199860 145024 199912
rect 145236 199860 145242 199912
rect 145294 199860 145300 199912
rect 145696 199860 145702 199912
rect 145754 199860 145760 199912
rect 145788 199860 145794 199912
rect 145846 199860 145852 199912
rect 145880 199860 145886 199912
rect 145938 199860 145944 199912
rect 145972 199860 145978 199912
rect 146030 199860 146036 199912
rect 146064 199860 146070 199912
rect 146122 199860 146128 199912
rect 144702 199832 144730 199860
rect 144702 199804 144960 199832
rect 144236 199600 144362 199628
rect 144236 199588 144242 199600
rect 144546 199588 144552 199640
rect 144604 199588 144610 199640
rect 142982 199520 142988 199572
rect 143040 199520 143046 199572
rect 144932 199504 144960 199804
rect 145254 199696 145282 199860
rect 145512 199792 145518 199844
rect 145570 199792 145576 199844
rect 145604 199792 145610 199844
rect 145662 199792 145668 199844
rect 145530 199708 145558 199792
rect 145254 199668 145328 199696
rect 145300 199640 145328 199668
rect 145466 199656 145472 199708
rect 145524 199668 145558 199708
rect 145524 199656 145530 199668
rect 145622 199640 145650 199792
rect 145282 199588 145288 199640
rect 145340 199588 145346 199640
rect 145558 199588 145564 199640
rect 145616 199600 145650 199640
rect 145616 199588 145622 199600
rect 145714 199572 145742 199860
rect 145806 199640 145834 199860
rect 145898 199696 145926 199860
rect 146082 199776 146110 199860
rect 146082 199736 146116 199776
rect 146110 199724 146116 199736
rect 146168 199724 146174 199776
rect 145898 199668 145972 199696
rect 145944 199640 145972 199668
rect 146018 199656 146024 199708
rect 146076 199696 146082 199708
rect 146220 199696 146248 199940
rect 147370 199912 147398 200212
rect 146340 199860 146346 199912
rect 146398 199860 146404 199912
rect 146708 199860 146714 199912
rect 146766 199860 146772 199912
rect 147168 199900 147174 199912
rect 147140 199860 147174 199900
rect 147226 199860 147232 199912
rect 147260 199860 147266 199912
rect 147318 199860 147324 199912
rect 147352 199860 147358 199912
rect 147410 199860 147416 199912
rect 147720 199860 147726 199912
rect 147778 199860 147784 199912
rect 148088 199860 148094 199912
rect 148146 199860 148152 199912
rect 148272 199860 148278 199912
rect 148330 199860 148336 199912
rect 148364 199860 148370 199912
rect 148422 199860 148428 199912
rect 146076 199668 146248 199696
rect 146076 199656 146082 199668
rect 145806 199600 145840 199640
rect 145834 199588 145840 199600
rect 145892 199588 145898 199640
rect 145926 199588 145932 199640
rect 145984 199588 145990 199640
rect 145650 199520 145656 199572
rect 145708 199532 145742 199572
rect 146358 199572 146386 199860
rect 146358 199532 146392 199572
rect 145708 199520 145714 199532
rect 146386 199520 146392 199532
rect 146444 199520 146450 199572
rect 146478 199520 146484 199572
rect 146536 199560 146542 199572
rect 146726 199560 146754 199860
rect 147140 199696 147168 199860
rect 147278 199832 147306 199860
rect 147232 199804 147306 199832
rect 147232 199776 147260 199804
rect 147214 199724 147220 199776
rect 147272 199724 147278 199776
rect 147738 199708 147766 199860
rect 147904 199792 147910 199844
rect 147962 199792 147968 199844
rect 147306 199696 147312 199708
rect 147140 199668 147312 199696
rect 147306 199656 147312 199668
rect 147364 199656 147370 199708
rect 147738 199668 147772 199708
rect 147766 199656 147772 199668
rect 147824 199656 147830 199708
rect 147922 199628 147950 199792
rect 148106 199708 148134 199860
rect 148290 199764 148318 199860
rect 148244 199736 148318 199764
rect 148244 199708 148272 199736
rect 148382 199708 148410 199860
rect 148042 199656 148048 199708
rect 148100 199668 148134 199708
rect 148100 199656 148106 199668
rect 148226 199656 148232 199708
rect 148284 199656 148290 199708
rect 148318 199656 148324 199708
rect 148376 199668 148410 199708
rect 148474 199696 148502 200348
rect 148566 199940 148686 199968
rect 148566 199912 148594 199940
rect 148548 199860 148554 199912
rect 148606 199860 148612 199912
rect 148548 199724 148554 199776
rect 148606 199764 148612 199776
rect 148658 199764 148686 199940
rect 149578 199912 149606 200416
rect 148916 199860 148922 199912
rect 148974 199860 148980 199912
rect 149284 199860 149290 199912
rect 149342 199860 149348 199912
rect 149468 199860 149474 199912
rect 149526 199860 149532 199912
rect 149560 199860 149566 199912
rect 149618 199860 149624 199912
rect 149836 199860 149842 199912
rect 149894 199860 149900 199912
rect 150020 199860 150026 199912
rect 150078 199860 150084 199912
rect 150480 199860 150486 199912
rect 150538 199860 150544 199912
rect 150572 199860 150578 199912
rect 150630 199860 150636 199912
rect 150664 199860 150670 199912
rect 150722 199860 150728 199912
rect 150848 199860 150854 199912
rect 150906 199860 150912 199912
rect 150940 199860 150946 199912
rect 150998 199860 151004 199912
rect 151032 199860 151038 199912
rect 151090 199860 151096 199912
rect 148934 199832 148962 199860
rect 148934 199804 149192 199832
rect 148606 199736 148686 199764
rect 148606 199724 148612 199736
rect 148474 199668 149008 199696
rect 148376 199656 148382 199668
rect 148980 199640 149008 199668
rect 148778 199628 148784 199640
rect 147922 199600 148784 199628
rect 148778 199588 148784 199600
rect 148836 199588 148842 199640
rect 148962 199588 148968 199640
rect 149020 199588 149026 199640
rect 149164 199572 149192 199804
rect 149302 199696 149330 199860
rect 149256 199668 149330 199696
rect 149486 199708 149514 199860
rect 149854 199776 149882 199860
rect 149854 199736 149888 199776
rect 149882 199724 149888 199736
rect 149940 199724 149946 199776
rect 149486 199668 149520 199708
rect 149256 199640 149284 199668
rect 149514 199656 149520 199668
rect 149572 199656 149578 199708
rect 150038 199696 150066 199860
rect 149716 199668 150066 199696
rect 149238 199588 149244 199640
rect 149296 199588 149302 199640
rect 149054 199560 149060 199572
rect 146536 199532 146754 199560
rect 148842 199532 149060 199560
rect 146536 199520 146542 199532
rect 142706 199492 142712 199504
rect 142586 199464 142712 199492
rect 142706 199452 142712 199464
rect 142764 199452 142770 199504
rect 144914 199452 144920 199504
rect 144972 199452 144978 199504
rect 136450 199384 136456 199436
rect 136508 199424 136514 199436
rect 148134 199424 148140 199436
rect 136508 199396 148140 199424
rect 136508 199384 136514 199396
rect 148134 199384 148140 199396
rect 148192 199384 148198 199436
rect 122742 199316 122748 199368
rect 122800 199356 122806 199368
rect 130010 199356 130016 199368
rect 122800 199328 130016 199356
rect 122800 199316 122806 199328
rect 130010 199316 130016 199328
rect 130068 199316 130074 199368
rect 133138 199316 133144 199368
rect 133196 199356 133202 199368
rect 133322 199356 133328 199368
rect 133196 199328 133328 199356
rect 133196 199316 133202 199328
rect 133322 199316 133328 199328
rect 133380 199316 133386 199368
rect 134610 199316 134616 199368
rect 134668 199328 134702 199368
rect 134668 199316 134674 199328
rect 139394 199316 139400 199368
rect 139452 199356 139458 199368
rect 139762 199356 139768 199368
rect 139452 199328 139768 199356
rect 139452 199316 139458 199328
rect 139762 199316 139768 199328
rect 139820 199316 139826 199368
rect 145098 199316 145104 199368
rect 145156 199356 145162 199368
rect 148842 199356 148870 199532
rect 149054 199520 149060 199532
rect 149112 199520 149118 199572
rect 149146 199520 149152 199572
rect 149204 199520 149210 199572
rect 149716 199560 149744 199668
rect 150296 199656 150302 199708
rect 150354 199656 150360 199708
rect 149790 199588 149796 199640
rect 149848 199628 149854 199640
rect 150314 199628 150342 199656
rect 149848 199600 150342 199628
rect 149848 199588 149854 199600
rect 150066 199560 150072 199572
rect 149716 199532 150072 199560
rect 150066 199520 150072 199532
rect 150124 199520 150130 199572
rect 150342 199520 150348 199572
rect 150400 199560 150406 199572
rect 150498 199560 150526 199860
rect 150400 199532 150526 199560
rect 150400 199520 150406 199532
rect 150590 199504 150618 199860
rect 148962 199452 148968 199504
rect 149020 199492 149026 199504
rect 149020 199452 149054 199492
rect 150526 199452 150532 199504
rect 150584 199464 150618 199504
rect 150584 199452 150590 199464
rect 145156 199328 148870 199356
rect 145156 199316 145162 199328
rect 122558 199248 122564 199300
rect 122616 199288 122622 199300
rect 145190 199288 145196 199300
rect 122616 199260 145196 199288
rect 122616 199248 122622 199260
rect 145190 199248 145196 199260
rect 145248 199248 145254 199300
rect 122466 199180 122472 199232
rect 122524 199220 122530 199232
rect 143442 199220 143448 199232
rect 122524 199192 143448 199220
rect 122524 199180 122530 199192
rect 143442 199180 143448 199192
rect 143500 199180 143506 199232
rect 149026 199220 149054 199452
rect 150682 199436 150710 199860
rect 150866 199832 150894 199860
rect 150820 199804 150894 199832
rect 150820 199640 150848 199804
rect 150958 199776 150986 199860
rect 150894 199724 150900 199776
rect 150952 199736 150986 199776
rect 150952 199724 150958 199736
rect 151050 199640 151078 199860
rect 151142 199696 151170 200484
rect 153442 200008 158990 200036
rect 151786 199940 153286 199968
rect 151676 199860 151682 199912
rect 151734 199860 151740 199912
rect 151142 199668 151584 199696
rect 151556 199640 151584 199668
rect 150802 199588 150808 199640
rect 150860 199588 150866 199640
rect 151050 199600 151084 199640
rect 151078 199588 151084 199600
rect 151136 199588 151142 199640
rect 151538 199588 151544 199640
rect 151596 199588 151602 199640
rect 150682 199396 150716 199436
rect 150710 199384 150716 199396
rect 150768 199384 150774 199436
rect 151694 199424 151722 199860
rect 150912 199396 151722 199424
rect 150912 199368 150940 199396
rect 150894 199316 150900 199368
rect 150952 199316 150958 199368
rect 151170 199316 151176 199368
rect 151228 199356 151234 199368
rect 151786 199356 151814 199940
rect 153258 199912 153286 199940
rect 153442 199912 153470 200008
rect 155282 199940 155678 199968
rect 151860 199860 151866 199912
rect 151918 199860 151924 199912
rect 151952 199860 151958 199912
rect 152010 199860 152016 199912
rect 152320 199860 152326 199912
rect 152378 199860 152384 199912
rect 152412 199860 152418 199912
rect 152470 199860 152476 199912
rect 152688 199860 152694 199912
rect 152746 199860 152752 199912
rect 152872 199860 152878 199912
rect 152930 199860 152936 199912
rect 153148 199860 153154 199912
rect 153206 199860 153212 199912
rect 153240 199860 153246 199912
rect 153298 199860 153304 199912
rect 153424 199860 153430 199912
rect 153482 199860 153488 199912
rect 153700 199860 153706 199912
rect 153758 199860 153764 199912
rect 153884 199860 153890 199912
rect 153942 199860 153948 199912
rect 154252 199860 154258 199912
rect 154310 199860 154316 199912
rect 154344 199860 154350 199912
rect 154402 199860 154408 199912
rect 155080 199860 155086 199912
rect 155138 199900 155144 199912
rect 155138 199872 155218 199900
rect 155138 199860 155144 199872
rect 151878 199776 151906 199860
rect 151970 199832 151998 199860
rect 151970 199804 152044 199832
rect 151878 199736 151912 199776
rect 151906 199724 151912 199736
rect 151964 199724 151970 199776
rect 152016 199708 152044 199804
rect 151998 199656 152004 199708
rect 152056 199656 152062 199708
rect 151228 199328 151814 199356
rect 151228 199316 151234 199328
rect 151538 199248 151544 199300
rect 151596 199288 151602 199300
rect 152338 199288 152366 199860
rect 152430 199708 152458 199860
rect 152430 199668 152464 199708
rect 152458 199656 152464 199668
rect 152516 199656 152522 199708
rect 152706 199560 152734 199860
rect 152890 199708 152918 199860
rect 152964 199792 152970 199844
rect 153022 199832 153028 199844
rect 153022 199792 153056 199832
rect 153028 199708 153056 199792
rect 152890 199668 152924 199708
rect 152918 199656 152924 199668
rect 152976 199656 152982 199708
rect 153010 199656 153016 199708
rect 153068 199656 153074 199708
rect 152826 199560 152832 199572
rect 152706 199532 152832 199560
rect 152826 199520 152832 199532
rect 152884 199520 152890 199572
rect 153166 199560 153194 199860
rect 153718 199776 153746 199860
rect 153654 199724 153660 199776
rect 153712 199736 153746 199776
rect 153712 199724 153718 199736
rect 153902 199640 153930 199860
rect 154068 199792 154074 199844
rect 154126 199792 154132 199844
rect 154086 199640 154114 199792
rect 154270 199776 154298 199860
rect 154206 199724 154212 199776
rect 154264 199736 154298 199776
rect 154264 199724 154270 199736
rect 154362 199640 154390 199860
rect 153838 199588 153844 199640
rect 153896 199600 153930 199640
rect 153896 199588 153902 199600
rect 154022 199588 154028 199640
rect 154080 199600 154114 199640
rect 154080 199588 154086 199600
rect 154298 199588 154304 199640
rect 154356 199600 154390 199640
rect 154850 199628 154856 199640
rect 154684 199600 154856 199628
rect 154356 199588 154362 199600
rect 154684 199572 154712 199600
rect 154850 199588 154856 199600
rect 154908 199588 154914 199640
rect 155190 199628 155218 199872
rect 155282 199776 155310 199940
rect 155650 199912 155678 199940
rect 156248 199940 157518 199968
rect 156248 199912 156276 199940
rect 155356 199860 155362 199912
rect 155414 199900 155420 199912
rect 155414 199872 155494 199900
rect 155414 199860 155420 199872
rect 155282 199736 155316 199776
rect 155310 199724 155316 199736
rect 155368 199724 155374 199776
rect 155466 199696 155494 199872
rect 155540 199860 155546 199912
rect 155598 199860 155604 199912
rect 155632 199860 155638 199912
rect 155690 199860 155696 199912
rect 156000 199860 156006 199912
rect 156058 199860 156064 199912
rect 156092 199860 156098 199912
rect 156150 199860 156156 199912
rect 156184 199860 156190 199912
rect 156242 199872 156276 199912
rect 156242 199860 156248 199872
rect 156368 199860 156374 199912
rect 156426 199860 156432 199912
rect 156644 199860 156650 199912
rect 156702 199860 156708 199912
rect 157380 199860 157386 199912
rect 157438 199860 157444 199912
rect 155558 199776 155586 199860
rect 155558 199736 155592 199776
rect 155586 199724 155592 199736
rect 155644 199724 155650 199776
rect 156018 199764 156046 199860
rect 156110 199832 156138 199860
rect 156276 199832 156282 199844
rect 156110 199804 156184 199832
rect 156156 199776 156184 199804
rect 156248 199792 156282 199832
rect 156334 199792 156340 199844
rect 156018 199736 156092 199764
rect 156064 199708 156092 199736
rect 156138 199724 156144 199776
rect 156196 199724 156202 199776
rect 156248 199708 156276 199792
rect 156386 199708 156414 199860
rect 155466 199668 156000 199696
rect 155862 199628 155868 199640
rect 155190 199600 155868 199628
rect 155862 199588 155868 199600
rect 155920 199588 155926 199640
rect 153378 199560 153384 199572
rect 153166 199532 153384 199560
rect 153378 199520 153384 199532
rect 153436 199520 153442 199572
rect 154666 199520 154672 199572
rect 154724 199520 154730 199572
rect 155402 199520 155408 199572
rect 155460 199560 155466 199572
rect 155972 199560 156000 199668
rect 156046 199656 156052 199708
rect 156104 199656 156110 199708
rect 156230 199656 156236 199708
rect 156288 199656 156294 199708
rect 156322 199656 156328 199708
rect 156380 199668 156414 199708
rect 156380 199656 156386 199668
rect 155460 199532 156000 199560
rect 156662 199560 156690 199860
rect 157398 199776 157426 199860
rect 157380 199724 157386 199776
rect 157438 199724 157444 199776
rect 156662 199532 157380 199560
rect 155460 199520 155466 199532
rect 154850 199452 154856 199504
rect 154908 199492 154914 199504
rect 154908 199464 154988 199492
rect 154908 199452 154914 199464
rect 154482 199384 154488 199436
rect 154540 199424 154546 199436
rect 154540 199396 154896 199424
rect 154540 199384 154546 199396
rect 154868 199368 154896 199396
rect 154850 199316 154856 199368
rect 154908 199316 154914 199368
rect 154960 199356 154988 199464
rect 156874 199384 156880 199436
rect 156932 199424 156938 199436
rect 157150 199424 157156 199436
rect 156932 199396 157156 199424
rect 156932 199384 156938 199396
rect 157150 199384 157156 199396
rect 157208 199384 157214 199436
rect 157242 199356 157248 199368
rect 154960 199328 157248 199356
rect 157242 199316 157248 199328
rect 157300 199316 157306 199368
rect 151596 199260 152366 199288
rect 151596 199248 151602 199260
rect 154390 199248 154396 199300
rect 154448 199288 154454 199300
rect 154758 199288 154764 199300
rect 154448 199260 154764 199288
rect 154448 199248 154454 199260
rect 154758 199248 154764 199260
rect 154816 199248 154822 199300
rect 156966 199248 156972 199300
rect 157024 199288 157030 199300
rect 157352 199288 157380 199532
rect 157024 199260 157380 199288
rect 157490 199288 157518 199940
rect 157564 199860 157570 199912
rect 157622 199860 157628 199912
rect 157748 199860 157754 199912
rect 157806 199860 157812 199912
rect 157840 199860 157846 199912
rect 157898 199860 157904 199912
rect 157932 199860 157938 199912
rect 157990 199860 157996 199912
rect 158024 199860 158030 199912
rect 158082 199860 158088 199912
rect 158208 199860 158214 199912
rect 158266 199860 158272 199912
rect 158300 199860 158306 199912
rect 158358 199860 158364 199912
rect 158484 199860 158490 199912
rect 158542 199860 158548 199912
rect 158668 199900 158674 199912
rect 158640 199860 158674 199900
rect 158726 199860 158732 199912
rect 158760 199860 158766 199912
rect 158818 199860 158824 199912
rect 158852 199860 158858 199912
rect 158910 199860 158916 199912
rect 157582 199356 157610 199860
rect 157766 199832 157794 199860
rect 157720 199804 157794 199832
rect 157720 199640 157748 199804
rect 157858 199708 157886 199860
rect 157794 199656 157800 199708
rect 157852 199668 157886 199708
rect 157852 199656 157858 199668
rect 157702 199588 157708 199640
rect 157760 199588 157766 199640
rect 157950 199628 157978 199860
rect 157812 199600 157978 199628
rect 157812 199492 157840 199600
rect 157886 199520 157892 199572
rect 157944 199560 157950 199572
rect 158042 199560 158070 199860
rect 158226 199640 158254 199860
rect 158162 199588 158168 199640
rect 158220 199600 158254 199640
rect 158220 199588 158226 199600
rect 157944 199532 158070 199560
rect 158318 199572 158346 199860
rect 158502 199640 158530 199860
rect 158438 199588 158444 199640
rect 158496 199600 158530 199640
rect 158496 199588 158502 199600
rect 158318 199532 158352 199572
rect 157944 199520 157950 199532
rect 158346 199520 158352 199532
rect 158404 199520 158410 199572
rect 158640 199504 158668 199860
rect 158778 199832 158806 199860
rect 158732 199804 158806 199832
rect 158732 199776 158760 199804
rect 158870 199776 158898 199860
rect 158714 199724 158720 199776
rect 158772 199724 158778 199776
rect 158806 199724 158812 199776
rect 158864 199736 158898 199776
rect 158864 199724 158870 199736
rect 158962 199572 158990 200008
rect 159128 199860 159134 199912
rect 159186 199860 159192 199912
rect 159312 199860 159318 199912
rect 159370 199860 159376 199912
rect 158898 199520 158904 199572
rect 158956 199532 158990 199572
rect 159146 199572 159174 199860
rect 159330 199640 159358 199860
rect 159422 199832 159450 200552
rect 159514 200484 173894 200512
rect 159514 199912 159542 200484
rect 173866 200444 173894 200484
rect 178954 200444 178960 200456
rect 173866 200416 178960 200444
rect 178954 200404 178960 200416
rect 179012 200404 179018 200456
rect 179386 200444 179414 200552
rect 180242 200444 180248 200456
rect 179386 200416 180248 200444
rect 180242 200404 180248 200416
rect 180300 200404 180306 200456
rect 187878 200376 187884 200388
rect 162274 200348 187884 200376
rect 159606 199940 159818 199968
rect 159496 199860 159502 199912
rect 159554 199860 159560 199912
rect 159606 199832 159634 199940
rect 159790 199844 159818 199940
rect 159956 199860 159962 199912
rect 160014 199860 160020 199912
rect 160048 199860 160054 199912
rect 160106 199860 160112 199912
rect 160140 199860 160146 199912
rect 160198 199860 160204 199912
rect 160508 199860 160514 199912
rect 160566 199860 160572 199912
rect 160784 199900 160790 199912
rect 160756 199860 160790 199900
rect 160842 199860 160848 199912
rect 160876 199860 160882 199912
rect 160934 199860 160940 199912
rect 160968 199860 160974 199912
rect 161026 199860 161032 199912
rect 161060 199860 161066 199912
rect 161118 199860 161124 199912
rect 161336 199860 161342 199912
rect 161394 199860 161400 199912
rect 161428 199860 161434 199912
rect 161486 199860 161492 199912
rect 161704 199860 161710 199912
rect 161762 199860 161768 199912
rect 161980 199860 161986 199912
rect 162038 199860 162044 199912
rect 159422 199804 159634 199832
rect 159680 199792 159686 199844
rect 159738 199792 159744 199844
rect 159772 199792 159778 199844
rect 159830 199792 159836 199844
rect 159864 199792 159870 199844
rect 159922 199792 159928 199844
rect 159588 199724 159594 199776
rect 159646 199724 159652 199776
rect 159606 199640 159634 199724
rect 159698 199708 159726 199792
rect 159882 199708 159910 199792
rect 159974 199776 160002 199860
rect 159956 199724 159962 199776
rect 160014 199724 160020 199776
rect 159698 199668 159732 199708
rect 159726 199656 159732 199668
rect 159784 199656 159790 199708
rect 159818 199656 159824 199708
rect 159876 199668 159910 199708
rect 160066 199696 160094 199860
rect 160158 199776 160186 199860
rect 160158 199736 160192 199776
rect 160186 199724 160192 199736
rect 160244 199724 160250 199776
rect 160020 199668 160094 199696
rect 159876 199656 159882 199668
rect 159330 199600 159364 199640
rect 159358 199588 159364 199600
rect 159416 199588 159422 199640
rect 159542 199588 159548 199640
rect 159600 199600 159634 199640
rect 159600 199588 159606 199600
rect 160020 199572 160048 199668
rect 159146 199532 159180 199572
rect 158956 199520 158962 199532
rect 159174 199520 159180 199532
rect 159232 199520 159238 199572
rect 160002 199520 160008 199572
rect 160060 199520 160066 199572
rect 160094 199520 160100 199572
rect 160152 199560 160158 199572
rect 160526 199560 160554 199860
rect 160600 199792 160606 199844
rect 160658 199792 160664 199844
rect 160152 199532 160554 199560
rect 160152 199520 160158 199532
rect 160618 199504 160646 199792
rect 160756 199504 160784 199860
rect 160894 199832 160922 199860
rect 160848 199804 160922 199832
rect 160848 199776 160876 199804
rect 160986 199776 161014 199860
rect 160830 199724 160836 199776
rect 160888 199724 160894 199776
rect 160922 199724 160928 199776
rect 160980 199736 161014 199776
rect 160980 199724 160986 199736
rect 161078 199708 161106 199860
rect 161354 199832 161382 199860
rect 161014 199656 161020 199708
rect 161072 199668 161106 199708
rect 161308 199804 161382 199832
rect 161072 199656 161078 199668
rect 161308 199572 161336 199804
rect 161446 199708 161474 199860
rect 161520 199792 161526 199844
rect 161578 199792 161584 199844
rect 161382 199656 161388 199708
rect 161440 199668 161474 199708
rect 161440 199656 161446 199668
rect 161538 199640 161566 199792
rect 161474 199588 161480 199640
rect 161532 199600 161566 199640
rect 161532 199588 161538 199600
rect 161290 199520 161296 199572
rect 161348 199520 161354 199572
rect 161722 199560 161750 199860
rect 161998 199708 162026 199860
rect 161934 199656 161940 199708
rect 161992 199668 162026 199708
rect 161992 199656 161998 199668
rect 161842 199560 161848 199572
rect 161722 199532 161848 199560
rect 161842 199520 161848 199532
rect 161900 199520 161906 199572
rect 162274 199504 162302 200348
rect 187878 200336 187884 200348
rect 187936 200336 187942 200388
rect 192110 200308 192116 200320
rect 164114 200280 192116 200308
rect 162458 199940 163038 199968
rect 162458 199912 162486 199940
rect 162348 199860 162354 199912
rect 162406 199860 162412 199912
rect 162440 199860 162446 199912
rect 162498 199860 162504 199912
rect 162532 199860 162538 199912
rect 162590 199900 162596 199912
rect 162716 199900 162722 199912
rect 162590 199860 162624 199900
rect 162366 199572 162394 199860
rect 162596 199640 162624 199860
rect 162688 199860 162722 199900
rect 162774 199860 162780 199912
rect 162808 199860 162814 199912
rect 162866 199860 162872 199912
rect 162900 199860 162906 199912
rect 162958 199860 162964 199912
rect 162688 199776 162716 199860
rect 162826 199832 162854 199860
rect 162780 199804 162854 199832
rect 162780 199776 162808 199804
rect 162918 199776 162946 199860
rect 162670 199724 162676 199776
rect 162728 199724 162734 199776
rect 162762 199724 162768 199776
rect 162820 199724 162826 199776
rect 162854 199724 162860 199776
rect 162912 199736 162946 199776
rect 162912 199724 162918 199736
rect 162578 199588 162584 199640
rect 162636 199588 162642 199640
rect 162366 199532 162400 199572
rect 162394 199520 162400 199532
rect 162452 199520 162458 199572
rect 163010 199504 163038 199940
rect 163470 199940 163774 199968
rect 163176 199860 163182 199912
rect 163234 199860 163240 199912
rect 163268 199860 163274 199912
rect 163326 199860 163332 199912
rect 163194 199708 163222 199860
rect 163286 199764 163314 199860
rect 163286 199736 163360 199764
rect 163194 199668 163228 199708
rect 163222 199656 163228 199668
rect 163280 199656 163286 199708
rect 163332 199640 163360 199736
rect 163314 199588 163320 199640
rect 163372 199588 163378 199640
rect 163470 199628 163498 199940
rect 163746 199912 163774 199940
rect 163544 199860 163550 199912
rect 163602 199860 163608 199912
rect 163636 199860 163642 199912
rect 163694 199860 163700 199912
rect 163728 199860 163734 199912
rect 163786 199860 163792 199912
rect 164004 199860 164010 199912
rect 164062 199860 164068 199912
rect 163562 199708 163590 199860
rect 163654 199764 163682 199860
rect 163654 199736 163912 199764
rect 163562 199668 163596 199708
rect 163590 199656 163596 199668
rect 163648 199656 163654 199708
rect 163884 199640 163912 199736
rect 163682 199628 163688 199640
rect 163470 199600 163688 199628
rect 163682 199588 163688 199600
rect 163740 199588 163746 199640
rect 163866 199588 163872 199640
rect 163924 199588 163930 199640
rect 157978 199492 157984 199504
rect 157812 199464 157984 199492
rect 157978 199452 157984 199464
rect 158036 199452 158042 199504
rect 158622 199452 158628 199504
rect 158680 199452 158686 199504
rect 160554 199452 160560 199504
rect 160612 199464 160646 199504
rect 160612 199452 160618 199464
rect 160738 199452 160744 199504
rect 160796 199452 160802 199504
rect 162274 199464 162308 199504
rect 162302 199452 162308 199464
rect 162360 199452 162366 199504
rect 163010 199464 163044 199504
rect 163038 199452 163044 199464
rect 163096 199452 163102 199504
rect 163774 199452 163780 199504
rect 163832 199492 163838 199504
rect 164022 199492 164050 199860
rect 163832 199464 164050 199492
rect 163832 199452 163838 199464
rect 159266 199384 159272 199436
rect 159324 199424 159330 199436
rect 159634 199424 159640 199436
rect 159324 199396 159640 199424
rect 159324 199384 159330 199396
rect 159634 199384 159640 199396
rect 159692 199384 159698 199436
rect 161566 199384 161572 199436
rect 161624 199424 161630 199436
rect 161750 199424 161756 199436
rect 161624 199396 161756 199424
rect 161624 199384 161630 199396
rect 161750 199384 161756 199396
rect 161808 199384 161814 199436
rect 162670 199384 162676 199436
rect 162728 199424 162734 199436
rect 162854 199424 162860 199436
rect 162728 199396 162860 199424
rect 162728 199384 162734 199396
rect 162854 199384 162860 199396
rect 162912 199384 162918 199436
rect 164114 199356 164142 200280
rect 192110 200268 192116 200280
rect 192168 200268 192174 200320
rect 190730 200240 190736 200252
rect 164666 200212 190736 200240
rect 164188 199860 164194 199912
rect 164246 199860 164252 199912
rect 164206 199424 164234 199860
rect 164372 199792 164378 199844
rect 164430 199792 164436 199844
rect 164390 199560 164418 199792
rect 164510 199560 164516 199572
rect 164390 199532 164516 199560
rect 164510 199520 164516 199532
rect 164568 199520 164574 199572
rect 164666 199492 164694 200212
rect 190730 200200 190736 200212
rect 190788 200200 190794 200252
rect 186774 200172 186780 200184
rect 167702 200144 186780 200172
rect 167702 199968 167730 200144
rect 186774 200132 186780 200144
rect 186832 200132 186838 200184
rect 178494 200104 178500 200116
rect 173130 200076 178500 200104
rect 165862 199940 166396 199968
rect 165862 199912 165890 199940
rect 164740 199860 164746 199912
rect 164798 199860 164804 199912
rect 164924 199860 164930 199912
rect 164982 199860 164988 199912
rect 165752 199860 165758 199912
rect 165810 199860 165816 199912
rect 165844 199860 165850 199912
rect 165902 199860 165908 199912
rect 165936 199860 165942 199912
rect 165994 199860 166000 199912
rect 166120 199860 166126 199912
rect 166178 199860 166184 199912
rect 164758 199560 164786 199860
rect 164942 199708 164970 199860
rect 165476 199792 165482 199844
rect 165534 199792 165540 199844
rect 164878 199656 164884 199708
rect 164936 199668 164970 199708
rect 164936 199656 164942 199668
rect 165062 199588 165068 199640
rect 165120 199628 165126 199640
rect 165494 199628 165522 199792
rect 165770 199776 165798 199860
rect 165954 199776 165982 199860
rect 165770 199736 165804 199776
rect 165798 199724 165804 199736
rect 165856 199724 165862 199776
rect 165890 199724 165896 199776
rect 165948 199736 165982 199776
rect 165948 199724 165954 199736
rect 166138 199696 166166 199860
rect 165120 199600 165522 199628
rect 165632 199668 166166 199696
rect 165120 199588 165126 199600
rect 165430 199560 165436 199572
rect 164758 199532 165436 199560
rect 165430 199520 165436 199532
rect 165488 199520 165494 199572
rect 164786 199492 164792 199504
rect 164666 199464 164792 199492
rect 164786 199452 164792 199464
rect 164844 199452 164850 199504
rect 165632 199492 165660 199668
rect 166368 199572 166396 199940
rect 166644 199940 167730 199968
rect 168116 199940 168558 199968
rect 166488 199860 166494 199912
rect 166546 199860 166552 199912
rect 166506 199640 166534 199860
rect 166644 199640 166672 199940
rect 167040 199900 167046 199912
rect 166736 199872 166948 199900
rect 166736 199640 166764 199872
rect 166442 199588 166448 199640
rect 166500 199600 166534 199640
rect 166500 199588 166506 199600
rect 166626 199588 166632 199640
rect 166684 199588 166690 199640
rect 166718 199588 166724 199640
rect 166776 199588 166782 199640
rect 166920 199572 166948 199872
rect 167012 199860 167046 199900
rect 167098 199860 167104 199912
rect 167224 199860 167230 199912
rect 167282 199860 167288 199912
rect 167316 199860 167322 199912
rect 167374 199860 167380 199912
rect 167592 199860 167598 199912
rect 167650 199860 167656 199912
rect 167960 199860 167966 199912
rect 168018 199860 168024 199912
rect 167012 199640 167040 199860
rect 167242 199776 167270 199860
rect 167178 199724 167184 199776
rect 167236 199736 167270 199776
rect 167334 199776 167362 199860
rect 167334 199736 167368 199776
rect 167236 199724 167242 199736
rect 167362 199724 167368 199736
rect 167420 199724 167426 199776
rect 166994 199588 167000 199640
rect 167052 199588 167058 199640
rect 166350 199520 166356 199572
rect 166408 199520 166414 199572
rect 166902 199520 166908 199572
rect 166960 199520 166966 199572
rect 167610 199560 167638 199860
rect 167978 199640 168006 199860
rect 167978 199600 168012 199640
rect 168006 199588 168012 199600
rect 168064 199588 168070 199640
rect 167610 199532 167684 199560
rect 166074 199492 166080 199504
rect 165632 199464 166080 199492
rect 166074 199452 166080 199464
rect 166132 199452 166138 199504
rect 165614 199424 165620 199436
rect 164206 199396 165620 199424
rect 165614 199384 165620 199396
rect 165672 199384 165678 199436
rect 167656 199368 167684 199532
rect 168116 199492 168144 199940
rect 168530 199912 168558 199940
rect 171658 199940 172974 199968
rect 171658 199912 171686 199940
rect 168420 199860 168426 199912
rect 168478 199860 168484 199912
rect 168512 199860 168518 199912
rect 168570 199860 168576 199912
rect 168604 199860 168610 199912
rect 168662 199860 168668 199912
rect 168788 199900 168794 199912
rect 168760 199860 168794 199900
rect 168846 199860 168852 199912
rect 168880 199860 168886 199912
rect 168938 199860 168944 199912
rect 168972 199860 168978 199912
rect 169030 199860 169036 199912
rect 169156 199900 169162 199912
rect 169128 199860 169162 199900
rect 169214 199860 169220 199912
rect 169248 199860 169254 199912
rect 169306 199860 169312 199912
rect 169340 199860 169346 199912
rect 169398 199860 169404 199912
rect 170168 199860 170174 199912
rect 170226 199860 170232 199912
rect 170536 199900 170542 199912
rect 170508 199860 170542 199900
rect 170594 199860 170600 199912
rect 170628 199860 170634 199912
rect 170686 199860 170692 199912
rect 170720 199860 170726 199912
rect 170778 199860 170784 199912
rect 171272 199860 171278 199912
rect 171330 199860 171336 199912
rect 171640 199860 171646 199912
rect 171698 199860 171704 199912
rect 171732 199860 171738 199912
rect 171790 199860 171796 199912
rect 172008 199900 172014 199912
rect 171980 199860 172014 199900
rect 172066 199860 172072 199912
rect 172192 199860 172198 199912
rect 172250 199860 172256 199912
rect 172744 199900 172750 199912
rect 172394 199872 172750 199900
rect 168190 199520 168196 199572
rect 168248 199560 168254 199572
rect 168438 199560 168466 199860
rect 168622 199708 168650 199860
rect 168558 199656 168564 199708
rect 168616 199668 168650 199708
rect 168616 199656 168622 199668
rect 168248 199532 168466 199560
rect 168248 199520 168254 199532
rect 168466 199492 168472 199504
rect 168116 199464 168472 199492
rect 168466 199452 168472 199464
rect 168524 199452 168530 199504
rect 168760 199492 168788 199860
rect 168898 199832 168926 199860
rect 168852 199804 168926 199832
rect 168852 199708 168880 199804
rect 168990 199708 169018 199860
rect 168834 199656 168840 199708
rect 168892 199656 168898 199708
rect 168926 199656 168932 199708
rect 168984 199668 169018 199708
rect 168984 199656 168990 199668
rect 169128 199640 169156 199860
rect 169266 199832 169294 199860
rect 169220 199804 169294 199832
rect 169220 199708 169248 199804
rect 169358 199708 169386 199860
rect 169202 199656 169208 199708
rect 169260 199656 169266 199708
rect 169294 199656 169300 199708
rect 169352 199668 169386 199708
rect 169352 199656 169358 199668
rect 169110 199588 169116 199640
rect 169168 199588 169174 199640
rect 170186 199560 170214 199860
rect 170352 199792 170358 199844
rect 170410 199832 170416 199844
rect 170410 199792 170444 199832
rect 170416 199640 170444 199792
rect 170508 199640 170536 199860
rect 170646 199832 170674 199860
rect 170600 199804 170674 199832
rect 170600 199708 170628 199804
rect 170738 199708 170766 199860
rect 170582 199656 170588 199708
rect 170640 199656 170646 199708
rect 170674 199656 170680 199708
rect 170732 199668 170766 199708
rect 170732 199656 170738 199668
rect 170398 199588 170404 199640
rect 170456 199588 170462 199640
rect 170490 199588 170496 199640
rect 170548 199588 170554 199640
rect 170858 199560 170864 199572
rect 170186 199532 170864 199560
rect 170858 199520 170864 199532
rect 170916 199520 170922 199572
rect 171290 199504 171318 199860
rect 171750 199776 171778 199860
rect 171686 199724 171692 199776
rect 171744 199736 171778 199776
rect 171744 199724 171750 199736
rect 171980 199572 172008 199860
rect 171962 199520 171968 199572
rect 172020 199520 172026 199572
rect 172210 199560 172238 199860
rect 172394 199696 172422 199872
rect 172744 199860 172750 199872
rect 172802 199860 172808 199912
rect 172836 199860 172842 199912
rect 172894 199860 172900 199912
rect 172854 199832 172882 199860
rect 172072 199532 172238 199560
rect 172348 199668 172422 199696
rect 172716 199804 172882 199832
rect 172072 199504 172100 199532
rect 169570 199492 169576 199504
rect 168760 199464 169576 199492
rect 169570 199452 169576 199464
rect 169628 199452 169634 199504
rect 171290 199464 171324 199504
rect 171318 199452 171324 199464
rect 171376 199452 171382 199504
rect 172054 199452 172060 199504
rect 172112 199452 172118 199504
rect 170030 199384 170036 199436
rect 170088 199424 170094 199436
rect 171870 199424 171876 199436
rect 170088 199396 171876 199424
rect 170088 199384 170094 199396
rect 171870 199384 171876 199396
rect 171928 199384 171934 199436
rect 172348 199424 172376 199668
rect 172716 199560 172744 199804
rect 172946 199628 172974 199940
rect 173020 199860 173026 199912
rect 173078 199900 173084 199912
rect 173130 199900 173158 200076
rect 178494 200064 178500 200076
rect 178552 200064 178558 200116
rect 178126 200036 178132 200048
rect 174832 200008 178132 200036
rect 173078 199872 173158 199900
rect 173078 199860 173084 199872
rect 173296 199860 173302 199912
rect 173354 199860 173360 199912
rect 173572 199860 173578 199912
rect 173630 199860 173636 199912
rect 173848 199860 173854 199912
rect 173906 199860 173912 199912
rect 173940 199860 173946 199912
rect 173998 199860 174004 199912
rect 174584 199860 174590 199912
rect 174642 199860 174648 199912
rect 174676 199860 174682 199912
rect 174734 199860 174740 199912
rect 173314 199696 173342 199860
rect 173314 199668 173480 199696
rect 172946 199600 173388 199628
rect 172974 199560 172980 199572
rect 172716 199532 172980 199560
rect 172974 199520 172980 199532
rect 173032 199520 173038 199572
rect 172422 199452 172428 199504
rect 172480 199492 172486 199504
rect 172790 199492 172796 199504
rect 172480 199464 172796 199492
rect 172480 199452 172486 199464
rect 172790 199452 172796 199464
rect 172848 199452 172854 199504
rect 172882 199424 172888 199436
rect 172348 199396 172888 199424
rect 172882 199384 172888 199396
rect 172940 199384 172946 199436
rect 173360 199424 173388 199600
rect 173452 199504 173480 199668
rect 173590 199560 173618 199860
rect 173866 199696 173894 199860
rect 173958 199832 173986 199860
rect 173958 199804 174032 199832
rect 173866 199668 173940 199696
rect 173912 199572 173940 199668
rect 174004 199640 174032 199804
rect 174124 199792 174130 199844
rect 174182 199792 174188 199844
rect 174142 199640 174170 199792
rect 174602 199764 174630 199860
rect 174280 199736 174630 199764
rect 173986 199588 173992 199640
rect 174044 199588 174050 199640
rect 174142 199600 174176 199640
rect 174170 199588 174176 199600
rect 174228 199588 174234 199640
rect 173802 199560 173808 199572
rect 173590 199532 173808 199560
rect 173802 199520 173808 199532
rect 173860 199520 173866 199572
rect 173894 199520 173900 199572
rect 173952 199520 173958 199572
rect 173434 199452 173440 199504
rect 173492 199452 173498 199504
rect 173710 199452 173716 199504
rect 173768 199492 173774 199504
rect 174280 199492 174308 199736
rect 174694 199708 174722 199860
rect 174630 199656 174636 199708
rect 174688 199668 174722 199708
rect 174688 199656 174694 199668
rect 174832 199640 174860 200008
rect 178126 199996 178132 200008
rect 178184 199996 178190 200048
rect 177942 199968 177948 199980
rect 175154 199940 175458 199968
rect 175154 199912 175182 199940
rect 174952 199860 174958 199912
rect 175010 199860 175016 199912
rect 175136 199860 175142 199912
rect 175194 199860 175200 199912
rect 175320 199860 175326 199912
rect 175378 199860 175384 199912
rect 174970 199696 174998 199860
rect 174924 199668 174998 199696
rect 174814 199588 174820 199640
rect 174872 199588 174878 199640
rect 174924 199560 174952 199668
rect 175338 199640 175366 199860
rect 175274 199588 175280 199640
rect 175332 199600 175366 199640
rect 175430 199628 175458 199940
rect 175522 199940 177948 199968
rect 175522 199912 175550 199940
rect 177942 199928 177948 199940
rect 178000 199928 178006 199980
rect 175504 199860 175510 199912
rect 175562 199860 175568 199912
rect 176056 199860 176062 199912
rect 176114 199860 176120 199912
rect 176240 199860 176246 199912
rect 176298 199860 176304 199912
rect 176424 199860 176430 199912
rect 176482 199860 176488 199912
rect 176700 199860 176706 199912
rect 176758 199860 176764 199912
rect 176884 199900 176890 199912
rect 176856 199860 176890 199900
rect 176942 199860 176948 199912
rect 176976 199860 176982 199912
rect 177034 199860 177040 199912
rect 177068 199860 177074 199912
rect 177126 199860 177132 199912
rect 175430 199600 175596 199628
rect 175332 199588 175338 199600
rect 175090 199560 175096 199572
rect 174924 199532 175096 199560
rect 175090 199520 175096 199532
rect 175148 199520 175154 199572
rect 173768 199464 174308 199492
rect 173768 199452 173774 199464
rect 174998 199452 175004 199504
rect 175056 199492 175062 199504
rect 175568 199492 175596 199600
rect 175056 199464 175596 199492
rect 176074 199492 176102 199860
rect 176258 199640 176286 199860
rect 176194 199588 176200 199640
rect 176252 199600 176286 199640
rect 176442 199640 176470 199860
rect 176718 199708 176746 199860
rect 176654 199656 176660 199708
rect 176712 199668 176746 199708
rect 176712 199656 176718 199668
rect 176442 199600 176476 199640
rect 176252 199588 176258 199600
rect 176470 199588 176476 199600
rect 176528 199588 176534 199640
rect 176856 199572 176884 199860
rect 176994 199832 177022 199860
rect 176948 199804 177022 199832
rect 176948 199708 176976 199804
rect 177086 199776 177114 199860
rect 177022 199724 177028 199776
rect 177080 199736 177114 199776
rect 177080 199724 177086 199736
rect 176930 199656 176936 199708
rect 176988 199656 176994 199708
rect 176838 199520 176844 199572
rect 176896 199520 176902 199572
rect 177298 199520 177304 199572
rect 177356 199560 177362 199572
rect 188154 199560 188160 199572
rect 177356 199532 188160 199560
rect 177356 199520 177362 199532
rect 188154 199520 188160 199532
rect 188212 199520 188218 199572
rect 177666 199492 177672 199504
rect 176074 199464 177672 199492
rect 175056 199452 175062 199464
rect 177666 199452 177672 199464
rect 177724 199452 177730 199504
rect 182910 199452 182916 199504
rect 182968 199492 182974 199504
rect 190546 199492 190552 199504
rect 182968 199464 190552 199492
rect 182968 199452 182974 199464
rect 190546 199452 190552 199464
rect 190604 199452 190610 199504
rect 179322 199424 179328 199436
rect 173360 199396 179328 199424
rect 179322 199384 179328 199396
rect 179380 199384 179386 199436
rect 180886 199384 180892 199436
rect 180944 199424 180950 199436
rect 190638 199424 190644 199436
rect 180944 199396 190644 199424
rect 180944 199384 180950 199396
rect 190638 199384 190644 199396
rect 190696 199384 190702 199436
rect 157582 199328 164142 199356
rect 167638 199316 167644 199368
rect 167696 199316 167702 199368
rect 170306 199316 170312 199368
rect 170364 199356 170370 199368
rect 200390 199356 200396 199368
rect 170364 199328 200396 199356
rect 170364 199316 170370 199328
rect 200390 199316 200396 199328
rect 200448 199316 200454 199368
rect 164786 199288 164792 199300
rect 157490 199260 164792 199288
rect 157024 199248 157030 199260
rect 164786 199248 164792 199260
rect 164844 199248 164850 199300
rect 167362 199248 167368 199300
rect 167420 199288 167426 199300
rect 201678 199288 201684 199300
rect 167420 199260 201684 199288
rect 167420 199248 167426 199260
rect 201678 199248 201684 199260
rect 201736 199248 201742 199300
rect 155310 199220 155316 199232
rect 149026 199192 155316 199220
rect 155310 199180 155316 199192
rect 155368 199180 155374 199232
rect 160002 199180 160008 199232
rect 160060 199220 160066 199232
rect 170398 199220 170404 199232
rect 160060 199192 170404 199220
rect 160060 199180 160066 199192
rect 170398 199180 170404 199192
rect 170456 199180 170462 199232
rect 172146 199180 172152 199232
rect 172204 199220 172210 199232
rect 180150 199220 180156 199232
rect 172204 199192 180156 199220
rect 172204 199180 172210 199192
rect 180150 199180 180156 199192
rect 180208 199180 180214 199232
rect 180794 199180 180800 199232
rect 180852 199220 180858 199232
rect 189810 199220 189816 199232
rect 180852 199192 189816 199220
rect 180852 199180 180858 199192
rect 189810 199180 189816 199192
rect 189868 199180 189874 199232
rect 122374 199112 122380 199164
rect 122432 199152 122438 199164
rect 145650 199152 145656 199164
rect 122432 199124 145656 199152
rect 122432 199112 122438 199124
rect 145650 199112 145656 199124
rect 145708 199112 145714 199164
rect 155862 199112 155868 199164
rect 155920 199152 155926 199164
rect 189074 199152 189080 199164
rect 155920 199124 189080 199152
rect 155920 199112 155926 199124
rect 189074 199112 189080 199124
rect 189132 199112 189138 199164
rect 121178 199044 121184 199096
rect 121236 199084 121242 199096
rect 132770 199084 132776 199096
rect 121236 199056 132776 199084
rect 121236 199044 121242 199056
rect 132770 199044 132776 199056
rect 132828 199044 132834 199096
rect 132954 199044 132960 199096
rect 133012 199084 133018 199096
rect 147582 199084 147588 199096
rect 133012 199056 147588 199084
rect 133012 199044 133018 199056
rect 147582 199044 147588 199056
rect 147640 199044 147646 199096
rect 150986 199044 150992 199096
rect 151044 199084 151050 199096
rect 158530 199084 158536 199096
rect 151044 199056 158536 199084
rect 151044 199044 151050 199056
rect 158530 199044 158536 199056
rect 158588 199044 158594 199096
rect 162302 199084 162308 199096
rect 158916 199056 162308 199084
rect 121270 198976 121276 199028
rect 121328 199016 121334 199028
rect 146570 199016 146576 199028
rect 121328 198988 146576 199016
rect 121328 198976 121334 198988
rect 146570 198976 146576 198988
rect 146628 198976 146634 199028
rect 153654 198976 153660 199028
rect 153712 199016 153718 199028
rect 158916 199016 158944 199056
rect 162302 199044 162308 199056
rect 162360 199044 162366 199096
rect 163130 199044 163136 199096
rect 163188 199084 163194 199096
rect 197538 199084 197544 199096
rect 163188 199056 197544 199084
rect 163188 199044 163194 199056
rect 197538 199044 197544 199056
rect 197596 199044 197602 199096
rect 153712 198988 158944 199016
rect 153712 198976 153718 198988
rect 158990 198976 158996 199028
rect 159048 199016 159054 199028
rect 193214 199016 193220 199028
rect 159048 198988 193220 199016
rect 159048 198976 159054 198988
rect 193214 198976 193220 198988
rect 193272 198976 193278 199028
rect 129550 198908 129556 198960
rect 129608 198948 129614 198960
rect 139026 198948 139032 198960
rect 129608 198920 139032 198948
rect 129608 198908 129614 198920
rect 139026 198908 139032 198920
rect 139084 198908 139090 198960
rect 139946 198908 139952 198960
rect 140004 198948 140010 198960
rect 144178 198948 144184 198960
rect 140004 198920 144184 198948
rect 140004 198908 140010 198920
rect 144178 198908 144184 198920
rect 144236 198908 144242 198960
rect 153930 198908 153936 198960
rect 153988 198948 153994 198960
rect 187786 198948 187792 198960
rect 153988 198920 187792 198948
rect 153988 198908 153994 198920
rect 187786 198908 187792 198920
rect 187844 198908 187850 198960
rect 129182 198840 129188 198892
rect 129240 198880 129246 198892
rect 147950 198880 147956 198892
rect 129240 198852 147956 198880
rect 129240 198840 129246 198852
rect 147950 198840 147956 198852
rect 148008 198840 148014 198892
rect 165982 198840 165988 198892
rect 166040 198880 166046 198892
rect 166718 198880 166724 198892
rect 166040 198852 166724 198880
rect 166040 198840 166046 198852
rect 166718 198840 166724 198852
rect 166776 198840 166782 198892
rect 170306 198880 170312 198892
rect 169680 198852 170312 198880
rect 126330 198772 126336 198824
rect 126388 198812 126394 198824
rect 144546 198812 144552 198824
rect 126388 198784 144552 198812
rect 126388 198772 126394 198784
rect 144546 198772 144552 198784
rect 144604 198772 144610 198824
rect 157242 198772 157248 198824
rect 157300 198772 157306 198824
rect 166074 198772 166080 198824
rect 166132 198812 166138 198824
rect 169680 198812 169708 198852
rect 170306 198840 170312 198852
rect 170364 198840 170370 198892
rect 170398 198840 170404 198892
rect 170456 198880 170462 198892
rect 172146 198880 172152 198892
rect 170456 198852 172152 198880
rect 170456 198840 170462 198852
rect 172146 198840 172152 198852
rect 172204 198840 172210 198892
rect 174446 198880 174452 198892
rect 172348 198852 174452 198880
rect 166132 198784 169708 198812
rect 166132 198772 166138 198784
rect 169754 198772 169760 198824
rect 169812 198812 169818 198824
rect 172348 198812 172376 198852
rect 174446 198840 174452 198852
rect 174504 198840 174510 198892
rect 174814 198880 174820 198892
rect 174556 198852 174820 198880
rect 169812 198784 172376 198812
rect 169812 198772 169818 198784
rect 172422 198772 172428 198824
rect 172480 198812 172486 198824
rect 172974 198812 172980 198824
rect 172480 198784 172980 198812
rect 172480 198772 172486 198784
rect 172974 198772 172980 198784
rect 173032 198772 173038 198824
rect 173250 198772 173256 198824
rect 173308 198812 173314 198824
rect 174556 198812 174584 198852
rect 174814 198840 174820 198852
rect 174872 198840 174878 198892
rect 175458 198840 175464 198892
rect 175516 198880 175522 198892
rect 180794 198880 180800 198892
rect 175516 198852 180800 198880
rect 175516 198840 175522 198852
rect 180794 198840 180800 198852
rect 180852 198840 180858 198892
rect 187510 198880 187516 198892
rect 180904 198852 187516 198880
rect 173308 198784 174584 198812
rect 173308 198772 173314 198784
rect 174630 198772 174636 198824
rect 174688 198812 174694 198824
rect 175642 198812 175648 198824
rect 174688 198784 175648 198812
rect 174688 198772 174694 198784
rect 175642 198772 175648 198784
rect 175700 198772 175706 198824
rect 175734 198772 175740 198824
rect 175792 198812 175798 198824
rect 176746 198812 176752 198824
rect 175792 198784 176752 198812
rect 175792 198772 175798 198784
rect 176746 198772 176752 198784
rect 176804 198772 176810 198824
rect 177942 198772 177948 198824
rect 178000 198812 178006 198824
rect 180904 198812 180932 198852
rect 187510 198840 187516 198852
rect 187568 198840 187574 198892
rect 178000 198784 180932 198812
rect 178000 198772 178006 198784
rect 183830 198772 183836 198824
rect 183888 198812 183894 198824
rect 189166 198812 189172 198824
rect 183888 198784 189172 198812
rect 183888 198772 183894 198784
rect 189166 198772 189172 198784
rect 189224 198772 189230 198824
rect 122650 198704 122656 198756
rect 122708 198744 122714 198756
rect 122708 198716 140774 198744
rect 122708 198704 122714 198716
rect 135070 198636 135076 198688
rect 135128 198676 135134 198688
rect 135254 198676 135260 198688
rect 135128 198648 135260 198676
rect 135128 198636 135134 198648
rect 135254 198636 135260 198648
rect 135312 198636 135318 198688
rect 140746 198676 140774 198716
rect 143718 198704 143724 198756
rect 143776 198744 143782 198756
rect 144086 198744 144092 198756
rect 143776 198716 144092 198744
rect 143776 198704 143782 198716
rect 144086 198704 144092 198716
rect 144144 198704 144150 198756
rect 157260 198744 157288 198772
rect 166626 198744 166632 198756
rect 157260 198716 166632 198744
rect 166626 198704 166632 198716
rect 166684 198704 166690 198756
rect 171410 198704 171416 198756
rect 171468 198744 171474 198756
rect 171468 198716 174584 198744
rect 171468 198704 171474 198716
rect 146202 198676 146208 198688
rect 140746 198648 146208 198676
rect 146202 198636 146208 198648
rect 146260 198636 146266 198688
rect 167178 198636 167184 198688
rect 167236 198676 167242 198688
rect 174170 198676 174176 198688
rect 167236 198648 174176 198676
rect 167236 198636 167242 198648
rect 174170 198636 174176 198648
rect 174228 198636 174234 198688
rect 174556 198676 174584 198716
rect 175918 198704 175924 198756
rect 175976 198744 175982 198756
rect 176470 198744 176476 198756
rect 175976 198716 176476 198744
rect 175976 198704 175982 198716
rect 176470 198704 176476 198716
rect 176528 198704 176534 198756
rect 177666 198704 177672 198756
rect 177724 198744 177730 198756
rect 201034 198744 201040 198756
rect 177724 198716 201040 198744
rect 177724 198704 177730 198716
rect 201034 198704 201040 198716
rect 201092 198704 201098 198756
rect 188338 198676 188344 198688
rect 174556 198648 188344 198676
rect 188338 198636 188344 198648
rect 188396 198636 188402 198688
rect 123110 198568 123116 198620
rect 123168 198608 123174 198620
rect 143626 198608 143632 198620
rect 123168 198580 143632 198608
rect 123168 198568 123174 198580
rect 143626 198568 143632 198580
rect 143684 198568 143690 198620
rect 148502 198568 148508 198620
rect 148560 198608 148566 198620
rect 149422 198608 149428 198620
rect 148560 198580 149428 198608
rect 148560 198568 148566 198580
rect 149422 198568 149428 198580
rect 149480 198568 149486 198620
rect 156782 198568 156788 198620
rect 156840 198608 156846 198620
rect 157150 198608 157156 198620
rect 156840 198580 157156 198608
rect 156840 198568 156846 198580
rect 157150 198568 157156 198580
rect 157208 198568 157214 198620
rect 167086 198568 167092 198620
rect 167144 198608 167150 198620
rect 170490 198608 170496 198620
rect 167144 198580 170496 198608
rect 167144 198568 167150 198580
rect 170490 198568 170496 198580
rect 170548 198568 170554 198620
rect 171870 198568 171876 198620
rect 171928 198608 171934 198620
rect 187050 198608 187056 198620
rect 171928 198580 187056 198608
rect 171928 198568 171934 198580
rect 187050 198568 187056 198580
rect 187108 198568 187114 198620
rect 108574 198500 108580 198552
rect 108632 198540 108638 198552
rect 128998 198540 129004 198552
rect 108632 198512 129004 198540
rect 108632 198500 108638 198512
rect 128998 198500 129004 198512
rect 129056 198500 129062 198552
rect 131758 198500 131764 198552
rect 131816 198540 131822 198552
rect 137554 198540 137560 198552
rect 131816 198512 137560 198540
rect 131816 198500 131822 198512
rect 137554 198500 137560 198512
rect 137612 198500 137618 198552
rect 137738 198500 137744 198552
rect 137796 198540 137802 198552
rect 138014 198540 138020 198552
rect 137796 198512 138020 198540
rect 137796 198500 137802 198512
rect 138014 198500 138020 198512
rect 138072 198500 138078 198552
rect 145650 198500 145656 198552
rect 145708 198540 145714 198552
rect 156690 198540 156696 198552
rect 145708 198512 156696 198540
rect 145708 198500 145714 198512
rect 156690 198500 156696 198512
rect 156748 198500 156754 198552
rect 171134 198500 171140 198552
rect 171192 198540 171198 198552
rect 186866 198540 186872 198552
rect 171192 198512 186872 198540
rect 171192 198500 171198 198512
rect 186866 198500 186872 198512
rect 186924 198500 186930 198552
rect 131850 198432 131856 198484
rect 131908 198472 131914 198484
rect 131908 198444 139624 198472
rect 131908 198432 131914 198444
rect 107102 198364 107108 198416
rect 107160 198404 107166 198416
rect 128538 198404 128544 198416
rect 107160 198376 128544 198404
rect 107160 198364 107166 198376
rect 128538 198364 128544 198376
rect 128596 198364 128602 198416
rect 130378 198364 130384 198416
rect 130436 198404 130442 198416
rect 138934 198404 138940 198416
rect 130436 198376 138940 198404
rect 130436 198364 130442 198376
rect 138934 198364 138940 198376
rect 138992 198364 138998 198416
rect 139596 198404 139624 198444
rect 141510 198432 141516 198484
rect 141568 198472 141574 198484
rect 142062 198472 142068 198484
rect 141568 198444 142068 198472
rect 141568 198432 141574 198444
rect 142062 198432 142068 198444
rect 142120 198432 142126 198484
rect 157794 198432 157800 198484
rect 157852 198472 157858 198484
rect 172422 198472 172428 198484
rect 157852 198444 172428 198472
rect 157852 198432 157858 198444
rect 172422 198432 172428 198444
rect 172480 198432 172486 198484
rect 174170 198432 174176 198484
rect 174228 198472 174234 198484
rect 178310 198472 178316 198484
rect 174228 198444 178316 198472
rect 174228 198432 174234 198444
rect 178310 198432 178316 198444
rect 178368 198432 178374 198484
rect 147674 198404 147680 198416
rect 139596 198376 147680 198404
rect 147674 198364 147680 198376
rect 147732 198364 147738 198416
rect 157058 198364 157064 198416
rect 157116 198404 157122 198416
rect 157426 198404 157432 198416
rect 157116 198376 157432 198404
rect 157116 198364 157122 198376
rect 157426 198364 157432 198376
rect 157484 198364 157490 198416
rect 158070 198364 158076 198416
rect 158128 198404 158134 198416
rect 173434 198404 173440 198416
rect 158128 198376 173440 198404
rect 158128 198364 158134 198376
rect 173434 198364 173440 198376
rect 173492 198364 173498 198416
rect 187970 198404 187976 198416
rect 173544 198376 187976 198404
rect 108666 198296 108672 198348
rect 108724 198336 108730 198348
rect 136450 198336 136456 198348
rect 108724 198308 136456 198336
rect 108724 198296 108730 198308
rect 136450 198296 136456 198308
rect 136508 198296 136514 198348
rect 136542 198296 136548 198348
rect 136600 198336 136606 198348
rect 145834 198336 145840 198348
rect 136600 198308 145840 198336
rect 136600 198296 136606 198308
rect 145834 198296 145840 198308
rect 145892 198296 145898 198348
rect 156414 198296 156420 198348
rect 156472 198336 156478 198348
rect 156472 198308 161474 198336
rect 156472 198296 156478 198308
rect 122098 198228 122104 198280
rect 122156 198268 122162 198280
rect 148502 198268 148508 198280
rect 122156 198240 148508 198268
rect 122156 198228 122162 198240
rect 148502 198228 148508 198240
rect 148560 198228 148566 198280
rect 151722 198228 151728 198280
rect 151780 198268 151786 198280
rect 158714 198268 158720 198280
rect 151780 198240 158720 198268
rect 151780 198228 151786 198240
rect 158714 198228 158720 198240
rect 158772 198228 158778 198280
rect 161446 198268 161474 198308
rect 170214 198296 170220 198348
rect 170272 198336 170278 198348
rect 173544 198336 173572 198376
rect 187970 198364 187976 198376
rect 188028 198364 188034 198416
rect 170272 198308 173572 198336
rect 170272 198296 170278 198308
rect 174446 198296 174452 198348
rect 174504 198336 174510 198348
rect 186958 198336 186964 198348
rect 174504 198308 186964 198336
rect 174504 198296 174510 198308
rect 186958 198296 186964 198308
rect 187016 198296 187022 198348
rect 161446 198240 167316 198268
rect 104434 198160 104440 198212
rect 104492 198200 104498 198212
rect 133230 198200 133236 198212
rect 104492 198172 133236 198200
rect 104492 198160 104498 198172
rect 133230 198160 133236 198172
rect 133288 198160 133294 198212
rect 138014 198160 138020 198212
rect 138072 198200 138078 198212
rect 139854 198200 139860 198212
rect 138072 198172 139860 198200
rect 138072 198160 138078 198172
rect 139854 198160 139860 198172
rect 139912 198160 139918 198212
rect 103054 198092 103060 198144
rect 103112 198132 103118 198144
rect 133966 198132 133972 198144
rect 103112 198104 133972 198132
rect 103112 198092 103118 198104
rect 133966 198092 133972 198104
rect 134024 198092 134030 198144
rect 146018 198132 146024 198144
rect 134076 198104 146024 198132
rect 103146 198024 103152 198076
rect 103204 198064 103210 198076
rect 128906 198064 128912 198076
rect 103204 198036 128912 198064
rect 103204 198024 103210 198036
rect 128906 198024 128912 198036
rect 128964 198024 128970 198076
rect 132770 198024 132776 198076
rect 132828 198064 132834 198076
rect 134076 198064 134104 198104
rect 146018 198092 146024 198104
rect 146076 198092 146082 198144
rect 167288 198132 167316 198240
rect 170766 198228 170772 198280
rect 170824 198268 170830 198280
rect 188062 198268 188068 198280
rect 170824 198240 188068 198268
rect 170824 198228 170830 198240
rect 188062 198228 188068 198240
rect 188120 198228 188126 198280
rect 170398 198160 170404 198212
rect 170456 198200 170462 198212
rect 188430 198200 188436 198212
rect 170456 198172 188436 198200
rect 170456 198160 170462 198172
rect 188430 198160 188436 198172
rect 188488 198160 188494 198212
rect 171042 198132 171048 198144
rect 164896 198104 167224 198132
rect 167288 198104 171048 198132
rect 132828 198036 134104 198064
rect 132828 198024 132834 198036
rect 140774 198024 140780 198076
rect 140832 198064 140838 198076
rect 141142 198064 141148 198076
rect 140832 198036 141148 198064
rect 140832 198024 140838 198036
rect 141142 198024 141148 198036
rect 141200 198024 141206 198076
rect 155954 198024 155960 198076
rect 156012 198064 156018 198076
rect 164896 198064 164924 198104
rect 156012 198036 164924 198064
rect 167196 198064 167224 198104
rect 171042 198092 171048 198104
rect 171100 198092 171106 198144
rect 172514 198092 172520 198144
rect 172572 198132 172578 198144
rect 172698 198132 172704 198144
rect 172572 198104 172704 198132
rect 172572 198092 172578 198104
rect 172698 198092 172704 198104
rect 172756 198092 172762 198144
rect 173894 198092 173900 198144
rect 173952 198132 173958 198144
rect 195330 198132 195336 198144
rect 173952 198104 195336 198132
rect 173952 198092 173958 198104
rect 195330 198092 195336 198104
rect 195388 198092 195394 198144
rect 171134 198064 171140 198076
rect 167196 198036 171140 198064
rect 156012 198024 156018 198036
rect 171134 198024 171140 198036
rect 171192 198024 171198 198076
rect 171318 198024 171324 198076
rect 171376 198064 171382 198076
rect 173250 198064 173256 198076
rect 171376 198036 173256 198064
rect 171376 198024 171382 198036
rect 173250 198024 173256 198036
rect 173308 198024 173314 198076
rect 198090 198064 198096 198076
rect 178006 198036 198096 198064
rect 102778 197956 102784 198008
rect 102836 197996 102842 198008
rect 126146 197996 126152 198008
rect 102836 197968 126152 197996
rect 102836 197956 102842 197968
rect 126146 197956 126152 197968
rect 126204 197956 126210 198008
rect 139486 197956 139492 198008
rect 139544 197996 139550 198008
rect 140498 197996 140504 198008
rect 139544 197968 140504 197996
rect 139544 197956 139550 197968
rect 140498 197956 140504 197968
rect 140556 197956 140562 198008
rect 165338 197956 165344 198008
rect 165396 197996 165402 198008
rect 174170 197996 174176 198008
rect 165396 197968 174176 197996
rect 165396 197956 165402 197968
rect 174170 197956 174176 197968
rect 174228 197956 174234 198008
rect 175642 197956 175648 198008
rect 175700 197996 175706 198008
rect 178006 197996 178034 198036
rect 198090 198024 198096 198036
rect 198148 198024 198154 198076
rect 175700 197968 178034 197996
rect 175700 197956 175706 197968
rect 178494 197956 178500 198008
rect 178552 197996 178558 198008
rect 199102 197996 199108 198008
rect 178552 197968 199108 197996
rect 178552 197956 178558 197968
rect 199102 197956 199108 197968
rect 199160 197956 199166 198008
rect 128262 197888 128268 197940
rect 128320 197928 128326 197940
rect 148042 197928 148048 197940
rect 128320 197900 148048 197928
rect 128320 197888 128326 197900
rect 148042 197888 148048 197900
rect 148100 197888 148106 197940
rect 155402 197888 155408 197940
rect 155460 197928 155466 197940
rect 171594 197928 171600 197940
rect 155460 197900 171600 197928
rect 155460 197888 155466 197900
rect 171594 197888 171600 197900
rect 171652 197888 171658 197940
rect 179322 197888 179328 197940
rect 179380 197928 179386 197940
rect 186682 197928 186688 197940
rect 179380 197900 186688 197928
rect 179380 197888 179386 197900
rect 186682 197888 186688 197900
rect 186740 197888 186746 197940
rect 132218 197820 132224 197872
rect 132276 197860 132282 197872
rect 151446 197860 151452 197872
rect 132276 197832 151452 197860
rect 132276 197820 132282 197832
rect 151446 197820 151452 197832
rect 151504 197820 151510 197872
rect 173802 197820 173808 197872
rect 173860 197860 173866 197872
rect 187418 197860 187424 197872
rect 173860 197832 187424 197860
rect 173860 197820 173866 197832
rect 187418 197820 187424 197832
rect 187476 197820 187482 197872
rect 126790 197752 126796 197804
rect 126848 197792 126854 197804
rect 145282 197792 145288 197804
rect 126848 197764 145288 197792
rect 126848 197752 126854 197764
rect 145282 197752 145288 197764
rect 145340 197752 145346 197804
rect 159634 197752 159640 197804
rect 159692 197792 159698 197804
rect 173710 197792 173716 197804
rect 159692 197764 173716 197792
rect 159692 197752 159698 197764
rect 173710 197752 173716 197764
rect 173768 197752 173774 197804
rect 126698 197684 126704 197736
rect 126756 197724 126762 197736
rect 146662 197724 146668 197736
rect 126756 197696 146668 197724
rect 126756 197684 126762 197696
rect 146662 197684 146668 197696
rect 146720 197684 146726 197736
rect 153378 197684 153384 197736
rect 153436 197724 153442 197736
rect 179046 197724 179052 197736
rect 153436 197696 179052 197724
rect 153436 197684 153442 197696
rect 179046 197684 179052 197696
rect 179104 197684 179110 197736
rect 123662 197616 123668 197668
rect 123720 197656 123726 197668
rect 145098 197656 145104 197668
rect 123720 197628 145104 197656
rect 123720 197616 123726 197628
rect 145098 197616 145104 197628
rect 145156 197616 145162 197668
rect 165430 197616 165436 197668
rect 165488 197656 165494 197668
rect 178954 197656 178960 197668
rect 165488 197628 178960 197656
rect 165488 197616 165494 197628
rect 178954 197616 178960 197628
rect 179012 197616 179018 197668
rect 132770 197548 132776 197600
rect 132828 197588 132834 197600
rect 145926 197588 145932 197600
rect 132828 197560 145932 197588
rect 132828 197548 132834 197560
rect 145926 197548 145932 197560
rect 145984 197548 145990 197600
rect 175274 197548 175280 197600
rect 175332 197588 175338 197600
rect 175550 197588 175556 197600
rect 175332 197560 175556 197588
rect 175332 197548 175338 197560
rect 175550 197548 175556 197560
rect 175608 197548 175614 197600
rect 134794 197480 134800 197532
rect 134852 197520 134858 197532
rect 135346 197520 135352 197532
rect 134852 197492 135352 197520
rect 134852 197480 134858 197492
rect 135346 197480 135352 197492
rect 135404 197480 135410 197532
rect 136634 197480 136640 197532
rect 136692 197520 136698 197532
rect 137186 197520 137192 197532
rect 136692 197492 137192 197520
rect 136692 197480 136698 197492
rect 137186 197480 137192 197492
rect 137244 197480 137250 197532
rect 161474 197480 161480 197532
rect 161532 197520 161538 197532
rect 161750 197520 161756 197532
rect 161532 197492 161756 197520
rect 161532 197480 161538 197492
rect 161750 197480 161756 197492
rect 161808 197480 161814 197532
rect 167730 197480 167736 197532
rect 167788 197520 167794 197532
rect 180610 197520 180616 197532
rect 167788 197492 180616 197520
rect 167788 197480 167794 197492
rect 180610 197480 180616 197492
rect 180668 197480 180674 197532
rect 162670 197412 162676 197464
rect 162728 197452 162734 197464
rect 163038 197452 163044 197464
rect 162728 197424 163044 197452
rect 162728 197412 162734 197424
rect 163038 197412 163044 197424
rect 163096 197412 163102 197464
rect 144546 197344 144552 197396
rect 144604 197384 144610 197396
rect 146938 197384 146944 197396
rect 144604 197356 146944 197384
rect 144604 197344 144610 197356
rect 146938 197344 146944 197356
rect 146996 197344 147002 197396
rect 147030 197344 147036 197396
rect 147088 197384 147094 197396
rect 147306 197384 147312 197396
rect 147088 197356 147312 197384
rect 147088 197344 147094 197356
rect 147306 197344 147312 197356
rect 147364 197344 147370 197396
rect 161474 197344 161480 197396
rect 161532 197384 161538 197396
rect 162026 197384 162032 197396
rect 161532 197356 162032 197384
rect 161532 197344 161538 197356
rect 162026 197344 162032 197356
rect 162084 197344 162090 197396
rect 162946 197344 162952 197396
rect 163004 197384 163010 197396
rect 163314 197384 163320 197396
rect 163004 197356 163320 197384
rect 163004 197344 163010 197356
rect 163314 197344 163320 197356
rect 163372 197344 163378 197396
rect 165706 197344 165712 197396
rect 165764 197384 165770 197396
rect 165982 197384 165988 197396
rect 165764 197356 165988 197384
rect 165764 197344 165770 197356
rect 165982 197344 165988 197356
rect 166040 197344 166046 197396
rect 171226 197344 171232 197396
rect 171284 197384 171290 197396
rect 171410 197384 171416 197396
rect 171284 197356 171416 197384
rect 171284 197344 171290 197356
rect 171410 197344 171416 197356
rect 171468 197344 171474 197396
rect 174078 197344 174084 197396
rect 174136 197384 174142 197396
rect 174354 197384 174360 197396
rect 174136 197356 174360 197384
rect 174136 197344 174142 197356
rect 174354 197344 174360 197356
rect 174412 197344 174418 197396
rect 175274 197344 175280 197396
rect 175332 197384 175338 197396
rect 175826 197384 175832 197396
rect 175332 197356 175832 197384
rect 175332 197344 175338 197356
rect 175826 197344 175832 197356
rect 175884 197344 175890 197396
rect 113818 197276 113824 197328
rect 113876 197316 113882 197328
rect 139210 197316 139216 197328
rect 113876 197288 139216 197316
rect 113876 197276 113882 197288
rect 139210 197276 139216 197288
rect 139268 197276 139274 197328
rect 160094 197276 160100 197328
rect 160152 197316 160158 197328
rect 161198 197316 161204 197328
rect 160152 197288 161204 197316
rect 160152 197276 160158 197288
rect 161198 197276 161204 197288
rect 161256 197276 161262 197328
rect 175366 197276 175372 197328
rect 175424 197316 175430 197328
rect 176562 197316 176568 197328
rect 175424 197288 176568 197316
rect 175424 197276 175430 197288
rect 176562 197276 176568 197288
rect 176620 197276 176626 197328
rect 176654 197276 176660 197328
rect 176712 197316 176718 197328
rect 179138 197316 179144 197328
rect 176712 197288 179144 197316
rect 176712 197276 176718 197288
rect 179138 197276 179144 197288
rect 179196 197276 179202 197328
rect 114186 197208 114192 197260
rect 114244 197248 114250 197260
rect 143166 197248 143172 197260
rect 114244 197220 143172 197248
rect 114244 197208 114250 197220
rect 143166 197208 143172 197220
rect 143224 197208 143230 197260
rect 163958 197208 163964 197260
rect 164016 197248 164022 197260
rect 194686 197248 194692 197260
rect 164016 197220 194692 197248
rect 164016 197208 164022 197220
rect 194686 197208 194692 197220
rect 194744 197208 194750 197260
rect 108390 197140 108396 197192
rect 108448 197180 108454 197192
rect 132954 197180 132960 197192
rect 108448 197152 132960 197180
rect 108448 197140 108454 197152
rect 132954 197140 132960 197152
rect 133012 197140 133018 197192
rect 138290 197180 138296 197192
rect 133064 197152 138296 197180
rect 114462 197072 114468 197124
rect 114520 197112 114526 197124
rect 132770 197112 132776 197124
rect 114520 197084 132776 197112
rect 114520 197072 114526 197084
rect 132770 197072 132776 197084
rect 132828 197072 132834 197124
rect 107194 197004 107200 197056
rect 107252 197044 107258 197056
rect 133064 197044 133092 197152
rect 138290 197140 138296 197152
rect 138348 197140 138354 197192
rect 162210 197140 162216 197192
rect 162268 197180 162274 197192
rect 194778 197180 194784 197192
rect 162268 197152 194784 197180
rect 162268 197140 162274 197152
rect 194778 197140 194784 197152
rect 194836 197140 194842 197192
rect 163498 197072 163504 197124
rect 163556 197112 163562 197124
rect 197354 197112 197360 197124
rect 163556 197084 197360 197112
rect 163556 197072 163562 197084
rect 197354 197072 197360 197084
rect 197412 197072 197418 197124
rect 107252 197016 133092 197044
rect 107252 197004 107258 197016
rect 133230 197004 133236 197056
rect 133288 197044 133294 197056
rect 143994 197044 144000 197056
rect 133288 197016 144000 197044
rect 133288 197004 133294 197016
rect 143994 197004 144000 197016
rect 144052 197004 144058 197056
rect 162854 197004 162860 197056
rect 162912 197044 162918 197056
rect 163774 197044 163780 197056
rect 162912 197016 163780 197044
rect 162912 197004 162918 197016
rect 163774 197004 163780 197016
rect 163832 197004 163838 197056
rect 168466 197004 168472 197056
rect 168524 197044 168530 197056
rect 168834 197044 168840 197056
rect 168524 197016 168840 197044
rect 168524 197004 168530 197016
rect 168834 197004 168840 197016
rect 168892 197004 168898 197056
rect 178954 197004 178960 197056
rect 179012 197044 179018 197056
rect 198826 197044 198832 197056
rect 179012 197016 198832 197044
rect 179012 197004 179018 197016
rect 198826 197004 198832 197016
rect 198884 197004 198890 197056
rect 111150 196936 111156 196988
rect 111208 196976 111214 196988
rect 142246 196976 142252 196988
rect 111208 196948 142252 196976
rect 111208 196936 111214 196948
rect 142246 196936 142252 196948
rect 142304 196936 142310 196988
rect 161934 196936 161940 196988
rect 161992 196976 161998 196988
rect 196066 196976 196072 196988
rect 161992 196948 196072 196976
rect 161992 196936 161998 196948
rect 196066 196936 196072 196948
rect 196124 196936 196130 196988
rect 117130 196868 117136 196920
rect 117188 196908 117194 196920
rect 149974 196908 149980 196920
rect 117188 196880 149980 196908
rect 117188 196868 117194 196880
rect 149974 196868 149980 196880
rect 150032 196868 150038 196920
rect 163866 196868 163872 196920
rect 163924 196908 163930 196920
rect 197446 196908 197452 196920
rect 163924 196880 197452 196908
rect 163924 196868 163930 196880
rect 197446 196868 197452 196880
rect 197504 196868 197510 196920
rect 110230 196800 110236 196852
rect 110288 196840 110294 196852
rect 144270 196840 144276 196852
rect 110288 196812 144276 196840
rect 110288 196800 110294 196812
rect 144270 196800 144276 196812
rect 144328 196800 144334 196852
rect 161382 196800 161388 196852
rect 161440 196840 161446 196852
rect 194594 196840 194600 196852
rect 161440 196812 194600 196840
rect 161440 196800 161446 196812
rect 194594 196800 194600 196812
rect 194652 196800 194658 196852
rect 105998 196732 106004 196784
rect 106056 196772 106062 196784
rect 139670 196772 139676 196784
rect 106056 196744 139676 196772
rect 106056 196732 106062 196744
rect 139670 196732 139676 196744
rect 139728 196732 139734 196784
rect 174170 196732 174176 196784
rect 174228 196772 174234 196784
rect 199010 196772 199016 196784
rect 174228 196744 199016 196772
rect 174228 196732 174234 196744
rect 199010 196732 199016 196744
rect 199068 196732 199074 196784
rect 110046 196664 110052 196716
rect 110104 196704 110110 196716
rect 133138 196704 133144 196716
rect 110104 196676 133144 196704
rect 110104 196664 110110 196676
rect 133138 196664 133144 196676
rect 133196 196664 133202 196716
rect 161658 196664 161664 196716
rect 161716 196704 161722 196716
rect 162394 196704 162400 196716
rect 161716 196676 162400 196704
rect 161716 196664 161722 196676
rect 162394 196664 162400 196676
rect 162452 196664 162458 196716
rect 164418 196664 164424 196716
rect 164476 196704 164482 196716
rect 198918 196704 198924 196716
rect 164476 196676 198924 196704
rect 164476 196664 164482 196676
rect 198918 196664 198924 196676
rect 198976 196664 198982 196716
rect 109954 196596 109960 196648
rect 110012 196636 110018 196648
rect 133230 196636 133236 196648
rect 110012 196608 133236 196636
rect 110012 196596 110018 196608
rect 133230 196596 133236 196608
rect 133288 196596 133294 196648
rect 161842 196596 161848 196648
rect 161900 196636 161906 196648
rect 196158 196636 196164 196648
rect 161900 196608 196164 196636
rect 161900 196596 161906 196608
rect 196158 196596 196164 196608
rect 196216 196596 196222 196648
rect 124858 196528 124864 196580
rect 124916 196568 124922 196580
rect 151078 196568 151084 196580
rect 124916 196540 151084 196568
rect 124916 196528 124922 196540
rect 151078 196528 151084 196540
rect 151136 196528 151142 196580
rect 123018 196460 123024 196512
rect 123076 196500 123082 196512
rect 143350 196500 143356 196512
rect 123076 196472 143356 196500
rect 123076 196460 123082 196472
rect 143350 196460 143356 196472
rect 143408 196460 143414 196512
rect 172422 196460 172428 196512
rect 172480 196500 172486 196512
rect 191926 196500 191932 196512
rect 172480 196472 191932 196500
rect 172480 196460 172486 196472
rect 191926 196460 191932 196472
rect 191984 196460 191990 196512
rect 129274 196392 129280 196444
rect 129332 196432 129338 196444
rect 145466 196432 145472 196444
rect 129332 196404 145472 196432
rect 129332 196392 129338 196404
rect 145466 196392 145472 196404
rect 145524 196392 145530 196444
rect 160002 196392 160008 196444
rect 160060 196432 160066 196444
rect 169938 196432 169944 196444
rect 160060 196404 169944 196432
rect 160060 196392 160066 196404
rect 169938 196392 169944 196404
rect 169996 196392 170002 196444
rect 173434 196392 173440 196444
rect 173492 196432 173498 196444
rect 191834 196432 191840 196444
rect 173492 196404 191840 196432
rect 173492 196392 173498 196404
rect 191834 196392 191840 196404
rect 191892 196392 191898 196444
rect 133138 196324 133144 196376
rect 133196 196364 133202 196376
rect 144638 196364 144644 196376
rect 133196 196336 144644 196364
rect 133196 196324 133202 196336
rect 144638 196324 144644 196336
rect 144696 196324 144702 196376
rect 164510 196324 164516 196376
rect 164568 196364 164574 196376
rect 180518 196364 180524 196376
rect 164568 196336 180524 196364
rect 164568 196324 164574 196336
rect 180518 196324 180524 196336
rect 180576 196324 180582 196376
rect 132954 196256 132960 196308
rect 133012 196296 133018 196308
rect 137738 196296 137744 196308
rect 133012 196268 137744 196296
rect 133012 196256 133018 196268
rect 137738 196256 137744 196268
rect 137796 196256 137802 196308
rect 160370 196256 160376 196308
rect 160428 196296 160434 196308
rect 169754 196296 169760 196308
rect 160428 196268 169760 196296
rect 160428 196256 160434 196268
rect 169754 196256 169760 196268
rect 169812 196256 169818 196308
rect 161106 196188 161112 196240
rect 161164 196228 161170 196240
rect 182818 196228 182824 196240
rect 161164 196200 182824 196228
rect 161164 196188 161170 196200
rect 182818 196188 182824 196200
rect 182876 196188 182882 196240
rect 160830 196120 160836 196172
rect 160888 196160 160894 196172
rect 183186 196160 183192 196172
rect 160888 196132 183192 196160
rect 160888 196120 160894 196132
rect 183186 196120 183192 196132
rect 183244 196120 183250 196172
rect 160370 196052 160376 196104
rect 160428 196092 160434 196104
rect 160922 196092 160928 196104
rect 160428 196064 160928 196092
rect 160428 196052 160434 196064
rect 160922 196052 160928 196064
rect 160980 196052 160986 196104
rect 171134 196052 171140 196104
rect 171192 196092 171198 196104
rect 171870 196092 171876 196104
rect 171192 196064 171876 196092
rect 171192 196052 171198 196064
rect 171870 196052 171876 196064
rect 171928 196052 171934 196104
rect 128722 195984 128728 196036
rect 128780 196024 128786 196036
rect 142430 196024 142436 196036
rect 128780 195996 142436 196024
rect 128780 195984 128786 195996
rect 142430 195984 142436 195996
rect 142488 195984 142494 196036
rect 146754 195984 146760 196036
rect 146812 196024 146818 196036
rect 147398 196024 147404 196036
rect 146812 195996 147404 196024
rect 146812 195984 146818 195996
rect 147398 195984 147404 195996
rect 147456 195984 147462 196036
rect 162762 195984 162768 196036
rect 162820 196024 162826 196036
rect 166994 196024 167000 196036
rect 162820 195996 167000 196024
rect 162820 195984 162826 195996
rect 166994 195984 167000 195996
rect 167052 195984 167058 196036
rect 112990 195916 112996 195968
rect 113048 195956 113054 195968
rect 142890 195956 142896 195968
rect 113048 195928 142896 195956
rect 113048 195916 113054 195928
rect 142890 195916 142896 195928
rect 142948 195916 142954 195968
rect 158898 195916 158904 195968
rect 158956 195956 158962 195968
rect 159818 195956 159824 195968
rect 158956 195928 159824 195956
rect 158956 195916 158962 195928
rect 159818 195916 159824 195928
rect 159876 195916 159882 195968
rect 171042 195916 171048 195968
rect 171100 195956 171106 195968
rect 190638 195956 190644 195968
rect 171100 195928 190644 195956
rect 171100 195916 171106 195928
rect 190638 195916 190644 195928
rect 190696 195916 190702 195968
rect 112806 195848 112812 195900
rect 112864 195888 112870 195900
rect 143074 195888 143080 195900
rect 112864 195860 143080 195888
rect 112864 195848 112870 195860
rect 143074 195848 143080 195860
rect 143132 195848 143138 195900
rect 156046 195848 156052 195900
rect 156104 195888 156110 195900
rect 157150 195888 157156 195900
rect 156104 195860 157156 195888
rect 156104 195848 156110 195860
rect 157150 195848 157156 195860
rect 157208 195848 157214 195900
rect 171870 195848 171876 195900
rect 171928 195888 171934 195900
rect 172146 195888 172152 195900
rect 171928 195860 172152 195888
rect 171928 195848 171934 195860
rect 172146 195848 172152 195860
rect 172204 195848 172210 195900
rect 172606 195848 172612 195900
rect 172664 195888 172670 195900
rect 172882 195888 172888 195900
rect 172664 195860 172888 195888
rect 172664 195848 172670 195860
rect 172882 195848 172888 195860
rect 172940 195848 172946 195900
rect 173710 195848 173716 195900
rect 173768 195888 173774 195900
rect 193306 195888 193312 195900
rect 173768 195860 193312 195888
rect 173768 195848 173774 195860
rect 193306 195848 193312 195860
rect 193364 195848 193370 195900
rect 108758 195780 108764 195832
rect 108816 195820 108822 195832
rect 140682 195820 140688 195832
rect 108816 195792 140688 195820
rect 108816 195780 108822 195792
rect 140682 195780 140688 195792
rect 140740 195780 140746 195832
rect 165614 195780 165620 195832
rect 165672 195820 165678 195832
rect 183278 195820 183284 195832
rect 165672 195792 183284 195820
rect 165672 195780 165678 195792
rect 183278 195780 183284 195792
rect 183336 195780 183342 195832
rect 108482 195712 108488 195764
rect 108540 195752 108546 195764
rect 140498 195752 140504 195764
rect 108540 195724 140504 195752
rect 108540 195712 108546 195724
rect 140498 195712 140504 195724
rect 140556 195712 140562 195764
rect 162670 195712 162676 195764
rect 162728 195752 162734 195764
rect 183002 195752 183008 195764
rect 162728 195724 183008 195752
rect 162728 195712 162734 195724
rect 183002 195712 183008 195724
rect 183060 195712 183066 195764
rect 100662 195644 100668 195696
rect 100720 195684 100726 195696
rect 133322 195684 133328 195696
rect 100720 195656 133328 195684
rect 100720 195644 100726 195656
rect 133322 195644 133328 195656
rect 133380 195644 133386 195696
rect 133966 195644 133972 195696
rect 134024 195684 134030 195696
rect 141050 195684 141056 195696
rect 134024 195656 141056 195684
rect 134024 195644 134030 195656
rect 141050 195644 141056 195656
rect 141108 195644 141114 195696
rect 159082 195644 159088 195696
rect 159140 195684 159146 195696
rect 159542 195684 159548 195696
rect 159140 195656 159548 195684
rect 159140 195644 159146 195656
rect 159542 195644 159548 195656
rect 159600 195644 159606 195696
rect 180242 195684 180248 195696
rect 171980 195656 180248 195684
rect 111518 195576 111524 195628
rect 111576 195616 111582 195628
rect 144086 195616 144092 195628
rect 111576 195588 144092 195616
rect 111576 195576 111582 195588
rect 144086 195576 144092 195588
rect 144144 195576 144150 195628
rect 154206 195576 154212 195628
rect 154264 195616 154270 195628
rect 154264 195588 161474 195616
rect 154264 195576 154270 195588
rect 112898 195508 112904 195560
rect 112956 195548 112962 195560
rect 145006 195548 145012 195560
rect 112956 195520 145012 195548
rect 112956 195508 112962 195520
rect 145006 195508 145012 195520
rect 145064 195508 145070 195560
rect 158622 195508 158628 195560
rect 158680 195548 158686 195560
rect 161446 195548 161474 195588
rect 171980 195548 172008 195656
rect 180242 195644 180248 195656
rect 180300 195644 180306 195696
rect 172054 195576 172060 195628
rect 172112 195616 172118 195628
rect 195146 195616 195152 195628
rect 172112 195588 195152 195616
rect 172112 195576 172118 195588
rect 195146 195576 195152 195588
rect 195204 195576 195210 195628
rect 158680 195520 159450 195548
rect 161446 195520 172008 195548
rect 158680 195508 158686 195520
rect 101674 195440 101680 195492
rect 101732 195480 101738 195492
rect 134150 195480 134156 195492
rect 101732 195452 134156 195480
rect 101732 195440 101738 195452
rect 134150 195440 134156 195452
rect 134208 195440 134214 195492
rect 159422 195480 159450 195520
rect 172146 195508 172152 195560
rect 172204 195548 172210 195560
rect 177298 195548 177304 195560
rect 172204 195520 177304 195548
rect 172204 195508 172210 195520
rect 177298 195508 177304 195520
rect 177356 195508 177362 195560
rect 190454 195480 190460 195492
rect 159422 195452 190460 195480
rect 190454 195440 190460 195452
rect 190512 195440 190518 195492
rect 105722 195372 105728 195424
rect 105780 195412 105786 195424
rect 139302 195412 139308 195424
rect 105780 195384 139308 195412
rect 105780 195372 105786 195384
rect 139302 195372 139308 195384
rect 139360 195372 139366 195424
rect 156598 195372 156604 195424
rect 156656 195412 156662 195424
rect 156656 195384 161474 195412
rect 156656 195372 156662 195384
rect 131850 195304 131856 195356
rect 131908 195344 131914 195356
rect 133966 195344 133972 195356
rect 131908 195316 133972 195344
rect 131908 195304 131914 195316
rect 133966 195304 133972 195316
rect 134024 195304 134030 195356
rect 134058 195304 134064 195356
rect 134116 195344 134122 195356
rect 134978 195344 134984 195356
rect 134116 195316 134984 195344
rect 134116 195304 134122 195316
rect 134978 195304 134984 195316
rect 135036 195304 135042 195356
rect 152918 195304 152924 195356
rect 152976 195344 152982 195356
rect 152976 195316 158576 195344
rect 152976 195304 152982 195316
rect 121362 195236 121368 195288
rect 121420 195276 121426 195288
rect 132034 195276 132040 195288
rect 121420 195248 132040 195276
rect 121420 195236 121426 195248
rect 132034 195236 132040 195248
rect 132092 195236 132098 195288
rect 134242 195236 134248 195288
rect 134300 195276 134306 195288
rect 134610 195276 134616 195288
rect 134300 195248 134616 195276
rect 134300 195236 134306 195248
rect 134610 195236 134616 195248
rect 134668 195236 134674 195288
rect 158070 195236 158076 195288
rect 158128 195276 158134 195288
rect 158438 195276 158444 195288
rect 158128 195248 158444 195276
rect 158128 195236 158134 195248
rect 158438 195236 158444 195248
rect 158496 195236 158502 195288
rect 158548 195276 158576 195316
rect 158806 195304 158812 195356
rect 158864 195344 158870 195356
rect 159358 195344 159364 195356
rect 158864 195316 159364 195344
rect 158864 195304 158870 195316
rect 159358 195304 159364 195316
rect 159416 195304 159422 195356
rect 161446 195344 161474 195384
rect 162578 195372 162584 195424
rect 162636 195412 162642 195424
rect 195974 195412 195980 195424
rect 162636 195384 195980 195412
rect 162636 195372 162642 195384
rect 195974 195372 195980 195384
rect 196032 195372 196038 195424
rect 190546 195344 190552 195356
rect 161446 195316 190552 195344
rect 190546 195304 190552 195316
rect 190604 195304 190610 195356
rect 186590 195276 186596 195288
rect 158548 195248 186596 195276
rect 186590 195236 186596 195248
rect 186648 195236 186654 195288
rect 122190 195168 122196 195220
rect 122248 195208 122254 195220
rect 148318 195208 148324 195220
rect 122248 195180 148324 195208
rect 122248 195168 122254 195180
rect 148318 195168 148324 195180
rect 148376 195168 148382 195220
rect 165614 195168 165620 195220
rect 165672 195208 165678 195220
rect 166718 195208 166724 195220
rect 165672 195180 166724 195208
rect 165672 195168 165678 195180
rect 166718 195168 166724 195180
rect 166776 195168 166782 195220
rect 169754 195168 169760 195220
rect 169812 195208 169818 195220
rect 172054 195208 172060 195220
rect 169812 195180 172060 195208
rect 169812 195168 169818 195180
rect 172054 195168 172060 195180
rect 172112 195168 172118 195220
rect 176838 195168 176844 195220
rect 176896 195208 176902 195220
rect 177206 195208 177212 195220
rect 176896 195180 177212 195208
rect 176896 195168 176902 195180
rect 177206 195168 177212 195180
rect 177264 195168 177270 195220
rect 177298 195168 177304 195220
rect 177356 195208 177362 195220
rect 189258 195208 189264 195220
rect 177356 195180 189264 195208
rect 177356 195168 177362 195180
rect 189258 195168 189264 195180
rect 189316 195168 189322 195220
rect 122282 195100 122288 195152
rect 122340 195140 122346 195152
rect 144822 195140 144828 195152
rect 122340 195112 144828 195140
rect 122340 195100 122346 195112
rect 144822 195100 144828 195112
rect 144880 195100 144886 195152
rect 164418 195100 164424 195152
rect 164476 195140 164482 195152
rect 165154 195140 165160 195152
rect 164476 195112 165160 195140
rect 164476 195100 164482 195112
rect 165154 195100 165160 195112
rect 165212 195100 165218 195152
rect 176746 195100 176752 195152
rect 176804 195140 176810 195152
rect 177574 195140 177580 195152
rect 176804 195112 177580 195140
rect 176804 195100 176810 195112
rect 177574 195100 177580 195112
rect 177632 195100 177638 195152
rect 126422 195032 126428 195084
rect 126480 195072 126486 195084
rect 144086 195072 144092 195084
rect 126480 195044 144092 195072
rect 126480 195032 126486 195044
rect 144086 195032 144092 195044
rect 144144 195032 144150 195084
rect 176654 195032 176660 195084
rect 176712 195072 176718 195084
rect 177666 195072 177672 195084
rect 176712 195044 177672 195072
rect 176712 195032 176718 195044
rect 177666 195032 177672 195044
rect 177724 195032 177730 195084
rect 121914 194964 121920 195016
rect 121972 195004 121978 195016
rect 156782 195004 156788 195016
rect 121972 194976 156788 195004
rect 121972 194964 121978 194976
rect 156782 194964 156788 194976
rect 156840 194964 156846 195016
rect 165706 194964 165712 195016
rect 165764 195004 165770 195016
rect 166442 195004 166448 195016
rect 165764 194976 166448 195004
rect 165764 194964 165770 194976
rect 166442 194964 166448 194976
rect 166500 194964 166506 195016
rect 171502 194964 171508 195016
rect 171560 195004 171566 195016
rect 189166 195004 189172 195016
rect 171560 194976 189172 195004
rect 171560 194964 171566 194976
rect 189166 194964 189172 194976
rect 189224 194964 189230 195016
rect 156138 194896 156144 194948
rect 156196 194936 156202 194948
rect 180426 194936 180432 194948
rect 156196 194908 180432 194936
rect 156196 194896 156202 194908
rect 180426 194896 180432 194908
rect 180484 194896 180490 194948
rect 106182 194488 106188 194540
rect 106240 194528 106246 194540
rect 136726 194528 136732 194540
rect 106240 194500 136732 194528
rect 106240 194488 106246 194500
rect 136726 194488 136732 194500
rect 136784 194488 136790 194540
rect 105906 194420 105912 194472
rect 105964 194460 105970 194472
rect 136910 194460 136916 194472
rect 105964 194432 136916 194460
rect 105964 194420 105970 194432
rect 136910 194420 136916 194432
rect 136968 194420 136974 194472
rect 103238 194352 103244 194404
rect 103296 194392 103302 194404
rect 135162 194392 135168 194404
rect 103296 194364 135168 194392
rect 103296 194352 103302 194364
rect 135162 194352 135168 194364
rect 135220 194352 135226 194404
rect 104526 194284 104532 194336
rect 104584 194324 104590 194336
rect 136082 194324 136088 194336
rect 104584 194296 136088 194324
rect 104584 194284 104590 194296
rect 136082 194284 136088 194296
rect 136140 194284 136146 194336
rect 104618 194216 104624 194268
rect 104676 194256 104682 194268
rect 135438 194256 135444 194268
rect 104676 194228 135444 194256
rect 104676 194216 104682 194228
rect 135438 194216 135444 194228
rect 135496 194216 135502 194268
rect 104158 194148 104164 194200
rect 104216 194188 104222 194200
rect 135898 194188 135904 194200
rect 104216 194160 135904 194188
rect 104216 194148 104222 194160
rect 135898 194148 135904 194160
rect 135956 194148 135962 194200
rect 102962 194080 102968 194132
rect 103020 194120 103026 194132
rect 134886 194120 134892 194132
rect 103020 194092 134892 194120
rect 103020 194080 103026 194092
rect 134886 194080 134892 194092
rect 134944 194080 134950 194132
rect 107010 194012 107016 194064
rect 107068 194052 107074 194064
rect 138014 194052 138020 194064
rect 107068 194024 138020 194052
rect 107068 194012 107074 194024
rect 138014 194012 138020 194024
rect 138072 194012 138078 194064
rect 103422 193944 103428 193996
rect 103480 193984 103486 193996
rect 136358 193984 136364 193996
rect 103480 193956 136364 193984
rect 103480 193944 103486 193956
rect 136358 193944 136364 193956
rect 136416 193944 136422 193996
rect 103330 193876 103336 193928
rect 103388 193916 103394 193928
rect 136634 193916 136640 193928
rect 103388 193888 136640 193916
rect 103388 193876 103394 193888
rect 136634 193876 136640 193888
rect 136692 193876 136698 193928
rect 168834 193876 168840 193928
rect 168892 193916 168898 193928
rect 203150 193916 203156 193928
rect 168892 193888 203156 193916
rect 168892 193876 168898 193888
rect 203150 193876 203156 193888
rect 203208 193876 203214 193928
rect 105814 193808 105820 193860
rect 105872 193848 105878 193860
rect 140222 193848 140228 193860
rect 105872 193820 140228 193848
rect 105872 193808 105878 193820
rect 140222 193808 140228 193820
rect 140280 193808 140286 193860
rect 168190 193808 168196 193860
rect 168248 193848 168254 193860
rect 201862 193848 201868 193860
rect 168248 193820 201868 193848
rect 168248 193808 168254 193820
rect 201862 193808 201868 193820
rect 201920 193808 201926 193860
rect 106918 193740 106924 193792
rect 106976 193780 106982 193792
rect 137462 193780 137468 193792
rect 106976 193752 137468 193780
rect 106976 193740 106982 193752
rect 137462 193740 137468 193752
rect 137520 193740 137526 193792
rect 104066 193672 104072 193724
rect 104124 193712 104130 193724
rect 128354 193712 128360 193724
rect 104124 193684 128360 193712
rect 104124 193672 104130 193684
rect 128354 193672 128360 193684
rect 128412 193672 128418 193724
rect 123386 193604 123392 193656
rect 123444 193644 123450 193656
rect 148226 193644 148232 193656
rect 123444 193616 148232 193644
rect 123444 193604 123450 193616
rect 148226 193604 148232 193616
rect 148284 193604 148290 193656
rect 145558 193196 145564 193248
rect 145616 193236 145622 193248
rect 149606 193236 149612 193248
rect 145616 193208 149612 193236
rect 145616 193196 145622 193208
rect 149606 193196 149612 193208
rect 149664 193196 149670 193248
rect 127710 193128 127716 193180
rect 127768 193168 127774 193180
rect 139486 193168 139492 193180
rect 127768 193140 139492 193168
rect 127768 193128 127774 193140
rect 139486 193128 139492 193140
rect 139544 193128 139550 193180
rect 163314 193128 163320 193180
rect 163372 193168 163378 193180
rect 179230 193168 179236 193180
rect 163372 193140 179236 193168
rect 163372 193128 163378 193140
rect 179230 193128 179236 193140
rect 179288 193128 179294 193180
rect 189718 193128 189724 193180
rect 189776 193168 189782 193180
rect 580166 193168 580172 193180
rect 189776 193140 580172 193168
rect 189776 193128 189782 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 114370 193060 114376 193112
rect 114428 193100 114434 193112
rect 143994 193100 144000 193112
rect 114428 193072 144000 193100
rect 114428 193060 114434 193072
rect 143994 193060 144000 193072
rect 144052 193060 144058 193112
rect 154390 193060 154396 193112
rect 154448 193100 154454 193112
rect 181530 193100 181536 193112
rect 154448 193072 181536 193100
rect 154448 193060 154454 193072
rect 181530 193060 181536 193072
rect 181588 193060 181594 193112
rect 115382 192992 115388 193044
rect 115440 193032 115446 193044
rect 146110 193032 146116 193044
rect 115440 193004 146116 193032
rect 115440 192992 115446 193004
rect 146110 192992 146116 193004
rect 146168 192992 146174 193044
rect 153286 192992 153292 193044
rect 153344 193032 153350 193044
rect 181622 193032 181628 193044
rect 153344 193004 181628 193032
rect 153344 192992 153350 193004
rect 181622 192992 181628 193004
rect 181680 192992 181686 193044
rect 101858 192924 101864 192976
rect 101916 192964 101922 192976
rect 134702 192964 134708 192976
rect 101916 192936 134708 192964
rect 101916 192924 101922 192936
rect 134702 192924 134708 192936
rect 134760 192924 134766 192976
rect 165430 192924 165436 192976
rect 165488 192964 165494 192976
rect 193858 192964 193864 192976
rect 165488 192936 193864 192964
rect 165488 192924 165494 192936
rect 193858 192924 193864 192936
rect 193916 192924 193922 192976
rect 116946 192856 116952 192908
rect 117004 192896 117010 192908
rect 149606 192896 149612 192908
rect 117004 192868 149612 192896
rect 117004 192856 117010 192868
rect 149606 192856 149612 192868
rect 149664 192856 149670 192908
rect 172882 192856 172888 192908
rect 172940 192896 172946 192908
rect 206094 192896 206100 192908
rect 172940 192868 206100 192896
rect 172940 192856 172946 192868
rect 206094 192856 206100 192868
rect 206152 192856 206158 192908
rect 111426 192788 111432 192840
rect 111484 192828 111490 192840
rect 143902 192828 143908 192840
rect 111484 192800 143908 192828
rect 111484 192788 111490 192800
rect 143902 192788 143908 192800
rect 143960 192788 143966 192840
rect 169386 192788 169392 192840
rect 169444 192828 169450 192840
rect 202874 192828 202880 192840
rect 169444 192800 202880 192828
rect 169444 192788 169450 192800
rect 202874 192788 202880 192800
rect 202932 192788 202938 192840
rect 109770 192720 109776 192772
rect 109828 192760 109834 192772
rect 142614 192760 142620 192772
rect 109828 192732 142620 192760
rect 109828 192720 109834 192732
rect 142614 192720 142620 192732
rect 142672 192720 142678 192772
rect 169018 192720 169024 192772
rect 169076 192760 169082 192772
rect 203058 192760 203064 192772
rect 169076 192732 203064 192760
rect 169076 192720 169082 192732
rect 203058 192720 203064 192732
rect 203116 192720 203122 192772
rect 117222 192652 117228 192704
rect 117280 192692 117286 192704
rect 150526 192692 150532 192704
rect 117280 192664 150532 192692
rect 117280 192652 117286 192664
rect 150526 192652 150532 192664
rect 150584 192652 150590 192704
rect 179690 192652 179696 192704
rect 179748 192692 179754 192704
rect 202414 192692 202420 192704
rect 179748 192664 202420 192692
rect 179748 192652 179754 192664
rect 202414 192652 202420 192664
rect 202472 192652 202478 192704
rect 108850 192584 108856 192636
rect 108908 192624 108914 192636
rect 142062 192624 142068 192636
rect 108908 192596 142068 192624
rect 108908 192584 108914 192596
rect 142062 192584 142068 192596
rect 142120 192584 142126 192636
rect 168742 192584 168748 192636
rect 168800 192624 168806 192636
rect 202966 192624 202972 192636
rect 168800 192596 202972 192624
rect 168800 192584 168806 192596
rect 202966 192584 202972 192596
rect 203024 192584 203030 192636
rect 109862 192516 109868 192568
rect 109920 192556 109926 192568
rect 144178 192556 144184 192568
rect 109920 192528 144184 192556
rect 109920 192516 109926 192528
rect 144178 192516 144184 192528
rect 144236 192516 144242 192568
rect 156322 192516 156328 192568
rect 156380 192556 156386 192568
rect 205634 192556 205640 192568
rect 156380 192528 205640 192556
rect 156380 192516 156386 192528
rect 205634 192516 205640 192528
rect 205692 192516 205698 192568
rect 112438 192448 112444 192500
rect 112496 192488 112502 192500
rect 144546 192488 144552 192500
rect 112496 192460 144552 192488
rect 112496 192448 112502 192460
rect 144546 192448 144552 192460
rect 144604 192448 144610 192500
rect 150710 192448 150716 192500
rect 150768 192488 150774 192500
rect 206186 192488 206192 192500
rect 150768 192460 206192 192488
rect 150768 192448 150774 192460
rect 206186 192448 206192 192460
rect 206244 192448 206250 192500
rect 114830 192380 114836 192432
rect 114888 192420 114894 192432
rect 144638 192420 144644 192432
rect 114888 192392 144644 192420
rect 114888 192380 114894 192392
rect 144638 192380 144644 192392
rect 144696 192380 144702 192432
rect 170490 192380 170496 192432
rect 170548 192420 170554 192432
rect 196802 192420 196808 192432
rect 170548 192392 196808 192420
rect 170548 192380 170554 192392
rect 196802 192380 196808 192392
rect 196860 192380 196866 192432
rect 127802 192312 127808 192364
rect 127860 192352 127866 192364
rect 139854 192352 139860 192364
rect 127860 192324 139860 192352
rect 127860 192312 127866 192324
rect 139854 192312 139860 192324
rect 139912 192312 139918 192364
rect 180610 192312 180616 192364
rect 180668 192352 180674 192364
rect 201586 192352 201592 192364
rect 180668 192324 201592 192352
rect 180668 192312 180674 192324
rect 201586 192312 201592 192324
rect 201644 192312 201650 192364
rect 130562 192244 130568 192296
rect 130620 192284 130626 192296
rect 140038 192284 140044 192296
rect 130620 192256 140044 192284
rect 130620 192244 130626 192256
rect 140038 192244 140044 192256
rect 140096 192244 140102 192296
rect 165798 192244 165804 192296
rect 165856 192284 165862 192296
rect 178954 192284 178960 192296
rect 165856 192256 178960 192284
rect 165856 192244 165862 192256
rect 178954 192244 178960 192256
rect 179012 192244 179018 192296
rect 149698 192176 149704 192228
rect 149756 192216 149762 192228
rect 151814 192216 151820 192228
rect 149756 192188 151820 192216
rect 149756 192176 149762 192188
rect 151814 192176 151820 192188
rect 151872 192176 151878 192228
rect 148962 191496 148968 191548
rect 149020 191536 149026 191548
rect 157610 191536 157616 191548
rect 149020 191508 157616 191536
rect 149020 191496 149026 191508
rect 157610 191496 157616 191508
rect 157668 191496 157674 191548
rect 115566 191428 115572 191480
rect 115624 191468 115630 191480
rect 139118 191468 139124 191480
rect 115624 191440 139124 191468
rect 115624 191428 115630 191440
rect 139118 191428 139124 191440
rect 139176 191428 139182 191480
rect 113082 191360 113088 191412
rect 113140 191400 113146 191412
rect 138934 191400 138940 191412
rect 113140 191372 138940 191400
rect 113140 191360 113146 191372
rect 138934 191360 138940 191372
rect 138992 191360 138998 191412
rect 111702 191292 111708 191344
rect 111760 191332 111766 191344
rect 138106 191332 138112 191344
rect 111760 191304 138112 191332
rect 111760 191292 111766 191304
rect 138106 191292 138112 191304
rect 138164 191292 138170 191344
rect 110322 191224 110328 191276
rect 110380 191264 110386 191276
rect 138382 191264 138388 191276
rect 110380 191236 138388 191264
rect 110380 191224 110386 191236
rect 138382 191224 138388 191236
rect 138440 191224 138446 191276
rect 150618 191224 150624 191276
rect 150676 191264 150682 191276
rect 151538 191264 151544 191276
rect 150676 191236 151544 191264
rect 150676 191224 150682 191236
rect 151538 191224 151544 191236
rect 151596 191224 151602 191276
rect 167270 191224 167276 191276
rect 167328 191264 167334 191276
rect 168282 191264 168288 191276
rect 167328 191236 168288 191264
rect 167328 191224 167334 191236
rect 168282 191224 168288 191236
rect 168340 191224 168346 191276
rect 104802 191156 104808 191208
rect 104860 191196 104866 191208
rect 137646 191196 137652 191208
rect 104860 191168 137652 191196
rect 104860 191156 104866 191168
rect 137646 191156 137652 191168
rect 137704 191156 137710 191208
rect 153286 191156 153292 191208
rect 153344 191196 153350 191208
rect 154298 191196 154304 191208
rect 153344 191168 154304 191196
rect 153344 191156 153350 191168
rect 154298 191156 154304 191168
rect 154356 191156 154362 191208
rect 169938 191156 169944 191208
rect 169996 191196 170002 191208
rect 170858 191196 170864 191208
rect 169996 191168 170864 191196
rect 169996 191156 170002 191168
rect 170858 191156 170864 191168
rect 170916 191156 170922 191208
rect 172514 191156 172520 191208
rect 172572 191196 172578 191208
rect 173342 191196 173348 191208
rect 172572 191168 173348 191196
rect 172572 191156 172578 191168
rect 173342 191156 173348 191168
rect 173400 191156 173406 191208
rect 174078 191156 174084 191208
rect 174136 191196 174142 191208
rect 174722 191196 174728 191208
rect 174136 191168 174728 191196
rect 174136 191156 174142 191168
rect 174722 191156 174728 191168
rect 174780 191156 174786 191208
rect 104342 191088 104348 191140
rect 104400 191128 104406 191140
rect 138658 191128 138664 191140
rect 104400 191100 138664 191128
rect 104400 191088 104406 191100
rect 138658 191088 138664 191100
rect 138716 191088 138722 191140
rect 169846 191088 169852 191140
rect 169904 191128 169910 191140
rect 170582 191128 170588 191140
rect 169904 191100 170588 191128
rect 169904 191088 169910 191100
rect 170582 191088 170588 191100
rect 170640 191088 170646 191140
rect 171318 191088 171324 191140
rect 171376 191128 171382 191140
rect 171962 191128 171968 191140
rect 171376 191100 171968 191128
rect 171376 191088 171382 191100
rect 171962 191088 171968 191100
rect 172020 191088 172026 191140
rect 172698 191088 172704 191140
rect 172756 191128 172762 191140
rect 173618 191128 173624 191140
rect 172756 191100 173624 191128
rect 172756 191088 172762 191100
rect 173618 191088 173624 191100
rect 173676 191088 173682 191140
rect 173986 191088 173992 191140
rect 174044 191128 174050 191140
rect 174446 191128 174452 191140
rect 174044 191100 174452 191128
rect 174044 191088 174050 191100
rect 174446 191088 174452 191100
rect 174504 191088 174510 191140
rect 175366 191088 175372 191140
rect 175424 191128 175430 191140
rect 176102 191128 176108 191140
rect 175424 191100 176108 191128
rect 175424 191088 175430 191100
rect 176102 191088 176108 191100
rect 176160 191088 176166 191140
rect 135622 191020 135628 191072
rect 135680 191060 135686 191072
rect 136174 191060 136180 191072
rect 135680 191032 136180 191060
rect 135680 191020 135686 191032
rect 136174 191020 136180 191032
rect 136232 191020 136238 191072
rect 142614 191020 142620 191072
rect 142672 191060 142678 191072
rect 143258 191060 143264 191072
rect 142672 191032 143264 191060
rect 142672 191020 142678 191032
rect 143258 191020 143264 191032
rect 143316 191020 143322 191072
rect 168466 191020 168472 191072
rect 168524 191060 168530 191072
rect 169202 191060 169208 191072
rect 168524 191032 169208 191060
rect 168524 191020 168530 191032
rect 169202 191020 169208 191032
rect 169260 191020 169266 191072
rect 170030 191020 170036 191072
rect 170088 191060 170094 191072
rect 170214 191060 170220 191072
rect 170088 191032 170220 191060
rect 170088 191020 170094 191032
rect 170214 191020 170220 191032
rect 170272 191020 170278 191072
rect 173894 191020 173900 191072
rect 173952 191060 173958 191072
rect 174998 191060 175004 191072
rect 173952 191032 175004 191060
rect 173952 191020 173958 191032
rect 174998 191020 175004 191032
rect 175056 191020 175062 191072
rect 110138 190136 110144 190188
rect 110196 190176 110202 190188
rect 141694 190176 141700 190188
rect 110196 190148 141700 190176
rect 110196 190136 110202 190148
rect 141694 190136 141700 190148
rect 141752 190136 141758 190188
rect 102870 190068 102876 190120
rect 102928 190108 102934 190120
rect 135530 190108 135536 190120
rect 102928 190080 135536 190108
rect 102928 190068 102934 190080
rect 135530 190068 135536 190080
rect 135588 190068 135594 190120
rect 101582 190000 101588 190052
rect 101640 190040 101646 190052
rect 134058 190040 134064 190052
rect 101640 190012 134064 190040
rect 101640 190000 101646 190012
rect 134058 190000 134064 190012
rect 134116 190000 134122 190052
rect 164326 190000 164332 190052
rect 164384 190040 164390 190052
rect 164602 190040 164608 190052
rect 164384 190012 164608 190040
rect 164384 190000 164390 190012
rect 164602 190000 164608 190012
rect 164660 190000 164666 190052
rect 108114 189932 108120 189984
rect 108172 189972 108178 189984
rect 141234 189972 141240 189984
rect 108172 189944 141240 189972
rect 108172 189932 108178 189944
rect 141234 189932 141240 189944
rect 141292 189932 141298 189984
rect 101950 189864 101956 189916
rect 102008 189904 102014 189916
rect 135806 189904 135812 189916
rect 102008 189876 135812 189904
rect 102008 189864 102014 189876
rect 135806 189864 135812 189876
rect 135864 189864 135870 189916
rect 171226 189864 171232 189916
rect 171284 189904 171290 189916
rect 172238 189904 172244 189916
rect 171284 189876 172244 189904
rect 171284 189864 171290 189876
rect 172238 189864 172244 189876
rect 172296 189864 172302 189916
rect 101766 189796 101772 189848
rect 101824 189836 101830 189848
rect 135346 189836 135352 189848
rect 101824 189808 135352 189836
rect 101824 189796 101830 189808
rect 135346 189796 135352 189808
rect 135404 189796 135410 189848
rect 106826 189728 106832 189780
rect 106884 189768 106890 189780
rect 141878 189768 141884 189780
rect 106884 189740 141884 189768
rect 106884 189728 106890 189740
rect 141878 189728 141884 189740
rect 141936 189728 141942 189780
rect 147582 189116 147588 189168
rect 147640 189156 147646 189168
rect 154758 189156 154764 189168
rect 147640 189128 154764 189156
rect 147640 189116 147646 189128
rect 154758 189116 154764 189128
rect 154816 189116 154822 189168
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 117866 189020 117872 189032
rect 3476 188992 117872 189020
rect 3476 188980 3482 188992
rect 117866 188980 117872 188992
rect 117924 188980 117930 189032
rect 154850 187552 154856 187604
rect 154908 187592 154914 187604
rect 155678 187592 155684 187604
rect 154908 187564 155684 187592
rect 154908 187552 154914 187564
rect 155678 187552 155684 187564
rect 155736 187552 155742 187604
rect 160554 186872 160560 186924
rect 160612 186912 160618 186924
rect 180058 186912 180064 186924
rect 160612 186884 180064 186912
rect 160612 186872 160618 186884
rect 180058 186872 180064 186884
rect 180116 186872 180122 186924
rect 148594 185784 148600 185836
rect 148652 185824 148658 185836
rect 154666 185824 154672 185836
rect 148652 185796 154672 185824
rect 148652 185784 148658 185796
rect 154666 185784 154672 185796
rect 154724 185784 154730 185836
rect 152550 185648 152556 185700
rect 152608 185688 152614 185700
rect 153010 185688 153016 185700
rect 152608 185660 153016 185688
rect 152608 185648 152614 185660
rect 153010 185648 153016 185660
rect 153068 185648 153074 185700
rect 154758 185580 154764 185632
rect 154816 185620 154822 185632
rect 155494 185620 155500 185632
rect 154816 185592 155500 185620
rect 154816 185580 154822 185592
rect 155494 185580 155500 185592
rect 155552 185580 155558 185632
rect 153378 185444 153384 185496
rect 153436 185484 153442 185496
rect 154114 185484 154120 185496
rect 153436 185456 154120 185484
rect 153436 185444 153442 185456
rect 154114 185444 154120 185456
rect 154172 185444 154178 185496
rect 160186 185376 160192 185428
rect 160244 185416 160250 185428
rect 160646 185416 160652 185428
rect 160244 185388 160652 185416
rect 160244 185376 160250 185388
rect 160646 185376 160652 185388
rect 160704 185376 160710 185428
rect 148042 184900 148048 184952
rect 148100 184940 148106 184952
rect 148870 184940 148876 184952
rect 148100 184912 148876 184940
rect 148100 184900 148106 184912
rect 148870 184900 148876 184912
rect 148928 184900 148934 184952
rect 145742 184696 145748 184748
rect 145800 184736 145806 184748
rect 156230 184736 156236 184748
rect 145800 184708 156236 184736
rect 145800 184696 145806 184708
rect 156230 184696 156236 184708
rect 156288 184696 156294 184748
rect 126606 183472 126612 183524
rect 126664 183512 126670 183524
rect 137922 183512 137928 183524
rect 126664 183484 137928 183512
rect 126664 183472 126670 183484
rect 137922 183472 137928 183484
rect 137980 183472 137986 183524
rect 149790 183200 149796 183252
rect 149848 183240 149854 183252
rect 151170 183240 151176 183252
rect 149848 183212 151176 183240
rect 149848 183200 149854 183212
rect 151170 183200 151176 183212
rect 151228 183200 151234 183252
rect 163130 182384 163136 182436
rect 163188 182424 163194 182436
rect 163682 182424 163688 182436
rect 163188 182396 163688 182424
rect 163188 182384 163194 182396
rect 163682 182384 163688 182396
rect 163740 182384 163746 182436
rect 188522 178032 188528 178084
rect 188580 178072 188586 178084
rect 580166 178072 580172 178084
rect 188580 178044 580172 178072
rect 188580 178032 188586 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 189718 165588 189724 165640
rect 189776 165628 189782 165640
rect 580166 165628 580172 165640
rect 189776 165600 580172 165628
rect 189776 165588 189782 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 193766 156612 193772 156664
rect 193824 156652 193830 156664
rect 193950 156652 193956 156664
rect 193824 156624 193956 156652
rect 193824 156612 193830 156624
rect 193950 156612 193956 156624
rect 194008 156612 194014 156664
rect 168558 155388 168564 155440
rect 168616 155428 168622 155440
rect 203334 155428 203340 155440
rect 168616 155400 203340 155428
rect 168616 155388 168622 155400
rect 203334 155388 203340 155400
rect 203392 155388 203398 155440
rect 168650 155320 168656 155372
rect 168708 155360 168714 155372
rect 203518 155360 203524 155372
rect 168708 155332 203524 155360
rect 168708 155320 168714 155332
rect 203518 155320 203524 155332
rect 203576 155320 203582 155372
rect 168466 155252 168472 155304
rect 168524 155292 168530 155304
rect 203426 155292 203432 155304
rect 168524 155264 203432 155292
rect 168524 155252 168530 155264
rect 203426 155252 203432 155264
rect 203484 155252 203490 155304
rect 167270 155184 167276 155236
rect 167328 155224 167334 155236
rect 202322 155224 202328 155236
rect 167328 155196 202328 155224
rect 167328 155184 167334 155196
rect 202322 155184 202328 155196
rect 202380 155184 202386 155236
rect 161750 153144 161756 153196
rect 161808 153184 161814 153196
rect 184658 153184 184664 153196
rect 161808 153156 184664 153184
rect 161808 153144 161814 153156
rect 184658 153144 184664 153156
rect 184716 153144 184722 153196
rect 160462 153076 160468 153128
rect 160520 153116 160526 153128
rect 184198 153116 184204 153128
rect 160520 153088 184204 153116
rect 160520 153076 160526 153088
rect 184198 153076 184204 153088
rect 184256 153076 184262 153128
rect 161566 153008 161572 153060
rect 161624 153048 161630 153060
rect 185578 153048 185584 153060
rect 161624 153020 185584 153048
rect 161624 153008 161630 153020
rect 185578 153008 185584 153020
rect 185636 153008 185642 153060
rect 160370 152940 160376 152992
rect 160428 152980 160434 152992
rect 185762 152980 185768 152992
rect 160428 152952 185768 152980
rect 160428 152940 160434 152952
rect 185762 152940 185768 152952
rect 185820 152940 185826 152992
rect 163038 152872 163044 152924
rect 163096 152912 163102 152924
rect 198182 152912 198188 152924
rect 163096 152884 198188 152912
rect 163096 152872 163102 152884
rect 198182 152872 198188 152884
rect 198240 152872 198246 152924
rect 164510 152804 164516 152856
rect 164568 152844 164574 152856
rect 199562 152844 199568 152856
rect 164568 152816 199568 152844
rect 164568 152804 164574 152816
rect 199562 152804 199568 152816
rect 199620 152804 199626 152856
rect 165982 152736 165988 152788
rect 166040 152776 166046 152788
rect 200666 152776 200672 152788
rect 166040 152748 200672 152776
rect 166040 152736 166046 152748
rect 200666 152736 200672 152748
rect 200724 152736 200730 152788
rect 168374 152668 168380 152720
rect 168432 152708 168438 152720
rect 203794 152708 203800 152720
rect 168432 152680 203800 152708
rect 168432 152668 168438 152680
rect 203794 152668 203800 152680
rect 203852 152668 203858 152720
rect 167086 152600 167092 152652
rect 167144 152640 167150 152652
rect 202046 152640 202052 152652
rect 167144 152612 202052 152640
rect 167144 152600 167150 152612
rect 202046 152600 202052 152612
rect 202104 152600 202110 152652
rect 168282 152532 168288 152584
rect 168340 152572 168346 152584
rect 202230 152572 202236 152584
rect 168340 152544 202236 152572
rect 168340 152532 168346 152544
rect 202230 152532 202236 152544
rect 202288 152532 202294 152584
rect 162762 152464 162768 152516
rect 162820 152504 162826 152516
rect 202138 152504 202144 152516
rect 162820 152476 202144 152504
rect 162820 152464 162826 152476
rect 202138 152464 202144 152476
rect 202196 152464 202202 152516
rect 163222 152396 163228 152448
rect 163280 152436 163286 152448
rect 184290 152436 184296 152448
rect 163280 152408 184296 152436
rect 163280 152396 163286 152408
rect 184290 152396 184296 152408
rect 184348 152396 184354 152448
rect 160278 150356 160284 150408
rect 160336 150396 160342 150408
rect 185762 150396 185768 150408
rect 160336 150368 185768 150396
rect 160336 150356 160342 150368
rect 185762 150356 185768 150368
rect 185820 150356 185826 150408
rect 158990 150288 158996 150340
rect 159048 150328 159054 150340
rect 184382 150328 184388 150340
rect 159048 150300 184388 150328
rect 159048 150288 159054 150300
rect 184382 150288 184388 150300
rect 184440 150288 184446 150340
rect 158898 150220 158904 150272
rect 158956 150260 158962 150272
rect 184566 150260 184572 150272
rect 158956 150232 184572 150260
rect 158956 150220 158962 150232
rect 184566 150220 184572 150232
rect 184624 150220 184630 150272
rect 158806 150152 158812 150204
rect 158864 150192 158870 150204
rect 184750 150192 184756 150204
rect 158864 150164 184756 150192
rect 158864 150152 158870 150164
rect 184750 150152 184756 150164
rect 184808 150152 184814 150204
rect 176838 150084 176844 150136
rect 176896 150124 176902 150136
rect 203702 150124 203708 150136
rect 176896 150096 203708 150124
rect 176896 150084 176902 150096
rect 203702 150084 203708 150096
rect 203760 150084 203766 150136
rect 176930 150016 176936 150068
rect 176988 150056 176994 150068
rect 204346 150056 204352 150068
rect 176988 150028 204352 150056
rect 176988 150016 176994 150028
rect 204346 150016 204352 150028
rect 204404 150016 204410 150068
rect 175642 149948 175648 150000
rect 175700 149988 175706 150000
rect 203610 149988 203616 150000
rect 175700 149960 203616 149988
rect 175700 149948 175706 149960
rect 203610 149948 203616 149960
rect 203668 149948 203674 150000
rect 175458 149880 175464 149932
rect 175516 149920 175522 149932
rect 204530 149920 204536 149932
rect 175516 149892 204536 149920
rect 175516 149880 175522 149892
rect 204530 149880 204536 149892
rect 204588 149880 204594 149932
rect 171594 149812 171600 149864
rect 171652 149852 171658 149864
rect 203242 149852 203248 149864
rect 171652 149824 203248 149852
rect 171652 149812 171658 149824
rect 203242 149812 203248 149824
rect 203300 149812 203306 149864
rect 152090 149744 152096 149796
rect 152148 149784 152154 149796
rect 204622 149784 204628 149796
rect 152148 149756 204628 149784
rect 152148 149744 152154 149756
rect 204622 149744 204628 149756
rect 204680 149744 204686 149796
rect 149238 149676 149244 149728
rect 149296 149716 149302 149728
rect 204438 149716 204444 149728
rect 149296 149688 204444 149716
rect 149296 149676 149302 149688
rect 204438 149676 204444 149688
rect 204496 149676 204502 149728
rect 159082 149608 159088 149660
rect 159140 149648 159146 149660
rect 184474 149648 184480 149660
rect 159140 149620 184480 149648
rect 159140 149608 159146 149620
rect 184474 149608 184480 149620
rect 184532 149608 184538 149660
rect 3418 149064 3424 149116
rect 3476 149104 3482 149116
rect 9582 149104 9588 149116
rect 3476 149076 9588 149104
rect 3476 149064 3482 149076
rect 9582 149064 9588 149076
rect 9640 149064 9646 149116
rect 115014 148996 115020 149048
rect 115072 149036 115078 149048
rect 142614 149036 142620 149048
rect 115072 149008 142620 149036
rect 115072 148996 115078 149008
rect 142614 148996 142620 149008
rect 142672 148996 142678 149048
rect 165614 148996 165620 149048
rect 165672 149036 165678 149048
rect 187142 149036 187148 149048
rect 165672 149008 187148 149036
rect 165672 148996 165678 149008
rect 187142 148996 187148 149008
rect 187200 148996 187206 149048
rect 113542 148928 113548 148980
rect 113600 148968 113606 148980
rect 143074 148968 143080 148980
rect 113600 148940 143080 148968
rect 113600 148928 113606 148940
rect 143074 148928 143080 148940
rect 143132 148928 143138 148980
rect 161474 148928 161480 148980
rect 161532 148968 161538 148980
rect 195422 148968 195428 148980
rect 161532 148940 195428 148968
rect 161532 148928 161538 148940
rect 195422 148928 195428 148940
rect 195480 148928 195486 148980
rect 125042 148860 125048 148912
rect 125100 148900 125106 148912
rect 153378 148900 153384 148912
rect 125100 148872 153384 148900
rect 125100 148860 125106 148872
rect 153378 148860 153384 148872
rect 153436 148860 153442 148912
rect 165890 148860 165896 148912
rect 165948 148900 165954 148912
rect 200942 148900 200948 148912
rect 165948 148872 200948 148900
rect 165948 148860 165954 148872
rect 200942 148860 200948 148872
rect 201000 148860 201006 148912
rect 120442 148792 120448 148844
rect 120500 148832 120506 148844
rect 149790 148832 149796 148844
rect 120500 148804 149796 148832
rect 120500 148792 120506 148804
rect 149790 148792 149796 148804
rect 149848 148792 149854 148844
rect 166902 148792 166908 148844
rect 166960 148832 166966 148844
rect 200850 148832 200856 148844
rect 166960 148804 200856 148832
rect 166960 148792 166966 148804
rect 200850 148792 200856 148804
rect 200908 148792 200914 148844
rect 108206 148724 108212 148776
rect 108264 148764 108270 148776
rect 138382 148764 138388 148776
rect 108264 148736 138388 148764
rect 108264 148724 108270 148736
rect 138382 148724 138388 148736
rect 138440 148724 138446 148776
rect 164418 148724 164424 148776
rect 164476 148764 164482 148776
rect 199654 148764 199660 148776
rect 164476 148736 199660 148764
rect 164476 148724 164482 148736
rect 199654 148724 199660 148736
rect 199712 148724 199718 148776
rect 122006 148656 122012 148708
rect 122064 148696 122070 148708
rect 153470 148696 153476 148708
rect 122064 148668 153476 148696
rect 122064 148656 122070 148668
rect 153470 148656 153476 148668
rect 153528 148656 153534 148708
rect 167822 148656 167828 148708
rect 167880 148696 167886 148708
rect 201954 148696 201960 148708
rect 167880 148668 201960 148696
rect 167880 148656 167886 148668
rect 201954 148656 201960 148668
rect 202012 148656 202018 148708
rect 100202 148588 100208 148640
rect 100260 148628 100266 148640
rect 133690 148628 133696 148640
rect 100260 148600 133696 148628
rect 100260 148588 100266 148600
rect 133690 148588 133696 148600
rect 133748 148588 133754 148640
rect 162946 148588 162952 148640
rect 163004 148628 163010 148640
rect 198458 148628 198464 148640
rect 163004 148600 198464 148628
rect 163004 148588 163010 148600
rect 198458 148588 198464 148600
rect 198516 148588 198522 148640
rect 100386 148520 100392 148572
rect 100444 148560 100450 148572
rect 134242 148560 134248 148572
rect 100444 148532 134248 148560
rect 100444 148520 100450 148532
rect 134242 148520 134248 148532
rect 134300 148520 134306 148572
rect 165706 148520 165712 148572
rect 165764 148560 165770 148572
rect 200758 148560 200764 148572
rect 165764 148532 200764 148560
rect 165764 148520 165770 148532
rect 200758 148520 200764 148532
rect 200816 148520 200822 148572
rect 100294 148452 100300 148504
rect 100352 148492 100358 148504
rect 134426 148492 134432 148504
rect 100352 148464 134432 148492
rect 100352 148452 100358 148464
rect 134426 148452 134432 148464
rect 134484 148452 134490 148504
rect 164326 148452 164332 148504
rect 164384 148492 164390 148504
rect 199470 148492 199476 148504
rect 164384 148464 199476 148492
rect 164384 148452 164390 148464
rect 199470 148452 199476 148464
rect 199528 148452 199534 148504
rect 105630 148384 105636 148436
rect 105688 148424 105694 148436
rect 139762 148424 139768 148436
rect 105688 148396 139768 148424
rect 105688 148384 105694 148396
rect 139762 148384 139768 148396
rect 139820 148384 139826 148436
rect 164234 148384 164240 148436
rect 164292 148424 164298 148436
rect 199378 148424 199384 148436
rect 164292 148396 199384 148424
rect 164292 148384 164298 148396
rect 199378 148384 199384 148396
rect 199436 148384 199442 148436
rect 9582 148316 9588 148368
rect 9640 148356 9646 148368
rect 180886 148356 180892 148368
rect 9640 148328 180892 148356
rect 9640 148316 9646 148328
rect 180886 148316 180892 148328
rect 180944 148356 180950 148368
rect 199286 148356 199292 148368
rect 180944 148328 199292 148356
rect 180944 148316 180950 148328
rect 199286 148316 199292 148328
rect 199344 148316 199350 148368
rect 121730 148248 121736 148300
rect 121788 148288 121794 148300
rect 148318 148288 148324 148300
rect 121788 148260 148324 148288
rect 121788 148248 121794 148260
rect 148318 148248 148324 148260
rect 148376 148248 148382 148300
rect 179230 148248 179236 148300
rect 179288 148288 179294 148300
rect 194134 148288 194140 148300
rect 179288 148260 194140 148288
rect 179288 148248 179294 148260
rect 194134 148248 194140 148260
rect 194192 148248 194198 148300
rect 114922 148180 114928 148232
rect 114980 148220 114986 148232
rect 140958 148220 140964 148232
rect 114980 148192 140964 148220
rect 114980 148180 114986 148192
rect 140958 148180 140964 148192
rect 141016 148180 141022 148232
rect 112254 148112 112260 148164
rect 112312 148152 112318 148164
rect 135622 148152 135628 148164
rect 112312 148124 135628 148152
rect 112312 148112 112318 148124
rect 135622 148112 135628 148124
rect 135680 148112 135686 148164
rect 179138 147568 179144 147620
rect 179196 147608 179202 147620
rect 196434 147608 196440 147620
rect 179196 147580 196440 147608
rect 179196 147568 179202 147580
rect 196434 147568 196440 147580
rect 196492 147568 196498 147620
rect 171502 147500 171508 147552
rect 171560 147540 171566 147552
rect 179230 147540 179236 147552
rect 171560 147512 179236 147540
rect 171560 147500 171566 147512
rect 179230 147500 179236 147512
rect 179288 147500 179294 147552
rect 179322 147500 179328 147552
rect 179380 147540 179386 147552
rect 196526 147540 196532 147552
rect 179380 147512 196532 147540
rect 179380 147500 179386 147512
rect 196526 147500 196532 147512
rect 196584 147500 196590 147552
rect 178402 147432 178408 147484
rect 178460 147472 178466 147484
rect 197906 147472 197912 147484
rect 178460 147444 197912 147472
rect 178460 147432 178466 147444
rect 197906 147432 197912 147444
rect 197964 147432 197970 147484
rect 170122 147364 170128 147416
rect 170180 147404 170186 147416
rect 192754 147404 192760 147416
rect 170180 147376 192760 147404
rect 170180 147364 170186 147376
rect 192754 147364 192760 147376
rect 192812 147364 192818 147416
rect 178218 147296 178224 147348
rect 178276 147336 178282 147348
rect 200574 147336 200580 147348
rect 178276 147308 200580 147336
rect 178276 147296 178282 147308
rect 200574 147296 200580 147308
rect 200632 147296 200638 147348
rect 117958 147228 117964 147280
rect 118016 147268 118022 147280
rect 127526 147268 127532 147280
rect 118016 147240 127532 147268
rect 118016 147228 118022 147240
rect 127526 147228 127532 147240
rect 127584 147228 127590 147280
rect 178678 147268 178684 147280
rect 161446 147240 178684 147268
rect 115198 147160 115204 147212
rect 115256 147200 115262 147212
rect 131850 147200 131856 147212
rect 115256 147172 131856 147200
rect 115256 147160 115262 147172
rect 131850 147160 131856 147172
rect 131908 147160 131914 147212
rect 110874 147092 110880 147144
rect 110932 147132 110938 147144
rect 128354 147132 128360 147144
rect 110932 147104 128360 147132
rect 110932 147092 110938 147104
rect 128354 147092 128360 147104
rect 128412 147092 128418 147144
rect 117682 147024 117688 147076
rect 117740 147064 117746 147076
rect 142522 147064 142528 147076
rect 117740 147036 142528 147064
rect 117740 147024 117746 147036
rect 142522 147024 142528 147036
rect 142580 147024 142586 147076
rect 110874 146956 110880 147008
rect 110932 146996 110938 147008
rect 137094 146996 137100 147008
rect 110932 146968 137100 146996
rect 110932 146956 110938 146968
rect 137094 146956 137100 146968
rect 137152 146956 137158 147008
rect 117590 146888 117596 146940
rect 117648 146928 117654 146940
rect 146478 146928 146484 146940
rect 117648 146900 146484 146928
rect 117648 146888 117654 146900
rect 146478 146888 146484 146900
rect 146536 146888 146542 146940
rect 148594 146888 148600 146940
rect 148652 146928 148658 146940
rect 161446 146928 161474 147240
rect 178678 147228 178684 147240
rect 178736 147228 178742 147280
rect 179230 147228 179236 147280
rect 179288 147268 179294 147280
rect 194042 147268 194048 147280
rect 179288 147240 194048 147268
rect 179288 147228 179294 147240
rect 194042 147228 194048 147240
rect 194100 147228 194106 147280
rect 172974 147160 172980 147212
rect 173032 147200 173038 147212
rect 178770 147200 178776 147212
rect 173032 147172 178776 147200
rect 173032 147160 173038 147172
rect 178770 147160 178776 147172
rect 178828 147160 178834 147212
rect 196986 147200 196992 147212
rect 178880 147172 196992 147200
rect 172606 147092 172612 147144
rect 172664 147132 172670 147144
rect 178880 147132 178908 147172
rect 196986 147160 196992 147172
rect 197044 147160 197050 147212
rect 172664 147104 178908 147132
rect 172664 147092 172670 147104
rect 179230 147092 179236 147144
rect 179288 147132 179294 147144
rect 195514 147132 195520 147144
rect 179288 147104 195520 147132
rect 179288 147092 179294 147104
rect 195514 147092 195520 147104
rect 195572 147092 195578 147144
rect 172882 147024 172888 147076
rect 172940 147064 172946 147076
rect 197078 147064 197084 147076
rect 172940 147036 197084 147064
rect 172940 147024 172946 147036
rect 197078 147024 197084 147036
rect 197136 147024 197142 147076
rect 178862 146956 178868 147008
rect 178920 146996 178926 147008
rect 179046 146996 179052 147008
rect 178920 146968 179052 146996
rect 178920 146956 178926 146968
rect 179046 146956 179052 146968
rect 179104 146956 179110 147008
rect 198274 146996 198280 147008
rect 179156 146968 198280 146996
rect 148652 146900 161474 146928
rect 148652 146888 148658 146900
rect 172790 146820 172796 146872
rect 172848 146860 172854 146872
rect 179156 146860 179184 146968
rect 198274 146956 198280 146968
rect 198332 146956 198338 147008
rect 196710 146928 196716 146940
rect 172848 146832 179184 146860
rect 179340 146900 196716 146928
rect 172848 146820 172854 146832
rect 171410 146752 171416 146804
rect 171468 146792 171474 146804
rect 179230 146792 179236 146804
rect 171468 146764 179236 146792
rect 171468 146752 171474 146764
rect 179230 146752 179236 146764
rect 179288 146752 179294 146804
rect 178034 146684 178040 146736
rect 178092 146724 178098 146736
rect 179340 146724 179368 146900
rect 196710 146888 196716 146900
rect 196768 146888 196774 146940
rect 180518 146820 180524 146872
rect 180576 146860 180582 146872
rect 192846 146860 192852 146872
rect 180576 146832 192852 146860
rect 180576 146820 180582 146832
rect 192846 146820 192852 146832
rect 192904 146820 192910 146872
rect 178092 146696 179368 146724
rect 178092 146684 178098 146696
rect 128354 146344 128360 146396
rect 128412 146384 128418 146396
rect 580442 146384 580448 146396
rect 128412 146356 580448 146384
rect 128412 146344 128418 146356
rect 580442 146344 580448 146356
rect 580500 146344 580506 146396
rect 127526 146276 127532 146328
rect 127584 146316 127590 146328
rect 580258 146316 580264 146328
rect 127584 146288 580264 146316
rect 127584 146276 127590 146288
rect 580258 146276 580264 146288
rect 580316 146276 580322 146328
rect 113450 146208 113456 146260
rect 113508 146248 113514 146260
rect 127802 146248 127808 146260
rect 113508 146220 127808 146248
rect 113508 146208 113514 146220
rect 127802 146208 127808 146220
rect 127860 146208 127866 146260
rect 179506 146208 179512 146260
rect 179564 146248 179570 146260
rect 195054 146248 195060 146260
rect 179564 146220 195060 146248
rect 179564 146208 179570 146220
rect 195054 146208 195060 146220
rect 195112 146208 195118 146260
rect 115290 146140 115296 146192
rect 115348 146180 115354 146192
rect 128906 146180 128912 146192
rect 115348 146152 128912 146180
rect 115348 146140 115354 146152
rect 128906 146140 128912 146152
rect 128964 146140 128970 146192
rect 183830 146140 183836 146192
rect 183888 146180 183894 146192
rect 199194 146180 199200 146192
rect 183888 146152 199200 146180
rect 183888 146140 183894 146152
rect 199194 146140 199200 146152
rect 199252 146140 199258 146192
rect 112714 146072 112720 146124
rect 112772 146112 112778 146124
rect 129918 146112 129924 146124
rect 112772 146084 129924 146112
rect 112772 146072 112778 146084
rect 129918 146072 129924 146084
rect 129976 146072 129982 146124
rect 178310 146072 178316 146124
rect 178368 146112 178374 146124
rect 193950 146112 193956 146124
rect 178368 146084 193956 146112
rect 178368 146072 178374 146084
rect 193950 146072 193956 146084
rect 194008 146072 194014 146124
rect 112530 146004 112536 146056
rect 112588 146044 112594 146056
rect 131298 146044 131304 146056
rect 112588 146016 131304 146044
rect 112588 146004 112594 146016
rect 131298 146004 131304 146016
rect 131356 146004 131362 146056
rect 178586 146004 178592 146056
rect 178644 146044 178650 146056
rect 195238 146044 195244 146056
rect 178644 146016 195244 146044
rect 178644 146004 178650 146016
rect 195238 146004 195244 146016
rect 195296 146004 195302 146056
rect 113726 145936 113732 145988
rect 113784 145976 113790 145988
rect 131574 145976 131580 145988
rect 113784 145948 131580 145976
rect 113784 145936 113790 145948
rect 131574 145936 131580 145948
rect 131632 145936 131638 145988
rect 175274 145936 175280 145988
rect 175332 145976 175338 145988
rect 195330 145976 195336 145988
rect 175332 145948 195336 145976
rect 175332 145936 175338 145948
rect 195330 145936 195336 145948
rect 195388 145936 195394 145988
rect 112530 145868 112536 145920
rect 112588 145908 112594 145920
rect 131758 145908 131764 145920
rect 112588 145880 131764 145908
rect 112588 145868 112594 145880
rect 131758 145868 131764 145880
rect 131816 145868 131822 145920
rect 172514 145868 172520 145920
rect 172572 145908 172578 145920
rect 195054 145908 195060 145920
rect 172572 145880 195060 145908
rect 172572 145868 172578 145880
rect 195054 145868 195060 145880
rect 195112 145868 195118 145920
rect 119062 145800 119068 145852
rect 119120 145840 119126 145852
rect 151446 145840 151452 145852
rect 119120 145812 151452 145840
rect 119120 145800 119126 145812
rect 151446 145800 151452 145812
rect 151504 145800 151510 145852
rect 173986 145800 173992 145852
rect 174044 145840 174050 145852
rect 197998 145840 198004 145852
rect 174044 145812 198004 145840
rect 174044 145800 174050 145812
rect 197998 145800 198004 145812
rect 198056 145800 198062 145852
rect 117498 145732 117504 145784
rect 117556 145772 117562 145784
rect 149698 145772 149704 145784
rect 117556 145744 149704 145772
rect 117556 145732 117562 145744
rect 149698 145732 149704 145744
rect 149756 145732 149762 145784
rect 160186 145732 160192 145784
rect 160244 145772 160250 145784
rect 192938 145772 192944 145784
rect 160244 145744 192944 145772
rect 160244 145732 160250 145744
rect 192938 145732 192944 145744
rect 192996 145732 193002 145784
rect 118970 145664 118976 145716
rect 119028 145704 119034 145716
rect 153010 145704 153016 145716
rect 119028 145676 153016 145704
rect 119028 145664 119034 145676
rect 153010 145664 153016 145676
rect 153068 145664 153074 145716
rect 160646 145664 160652 145716
rect 160704 145704 160710 145716
rect 193398 145704 193404 145716
rect 160704 145676 193404 145704
rect 160704 145664 160710 145676
rect 193398 145664 193404 145676
rect 193456 145664 193462 145716
rect 116210 145596 116216 145648
rect 116268 145636 116274 145648
rect 147858 145636 147864 145648
rect 116268 145608 147864 145636
rect 116268 145596 116274 145608
rect 147858 145596 147864 145608
rect 147916 145596 147922 145648
rect 148962 145596 148968 145648
rect 149020 145636 149026 145648
rect 189994 145636 190000 145648
rect 149020 145608 190000 145636
rect 149020 145596 149026 145608
rect 189994 145596 190000 145608
rect 190052 145596 190058 145648
rect 3510 145528 3516 145580
rect 3568 145568 3574 145580
rect 3568 145540 161474 145568
rect 3568 145528 3574 145540
rect 161446 145432 161474 145540
rect 183462 145528 183468 145580
rect 183520 145568 183526 145580
rect 200482 145568 200488 145580
rect 183520 145540 200488 145568
rect 183520 145528 183526 145540
rect 200482 145528 200488 145540
rect 200540 145528 200546 145580
rect 179414 145460 179420 145512
rect 179472 145500 179478 145512
rect 194870 145500 194876 145512
rect 179472 145472 194876 145500
rect 179472 145460 179478 145472
rect 194870 145460 194876 145472
rect 194928 145460 194934 145512
rect 179598 145432 179604 145444
rect 161446 145404 179604 145432
rect 179598 145392 179604 145404
rect 179656 145432 179662 145444
rect 192478 145432 192484 145444
rect 179656 145404 192484 145432
rect 179656 145392 179662 145404
rect 192478 145392 192484 145404
rect 192536 145392 192542 145444
rect 120534 144916 120540 144968
rect 120592 144956 120598 144968
rect 182266 144956 182272 144968
rect 120592 144928 182272 144956
rect 120592 144916 120598 144928
rect 182266 144916 182272 144928
rect 182324 144956 182330 144968
rect 183462 144956 183468 144968
rect 182324 144928 183468 144956
rect 182324 144916 182330 144928
rect 183462 144916 183468 144928
rect 183520 144916 183526 144968
rect 184658 144848 184664 144900
rect 184716 144888 184722 144900
rect 196894 144888 196900 144900
rect 184716 144860 196900 144888
rect 184716 144848 184722 144860
rect 196894 144848 196900 144860
rect 196952 144848 196958 144900
rect 172422 144780 172428 144832
rect 172480 144820 172486 144832
rect 190822 144820 190828 144832
rect 172480 144792 190828 144820
rect 172480 144780 172486 144792
rect 190822 144780 190828 144792
rect 190880 144780 190886 144832
rect 112714 144712 112720 144764
rect 112772 144752 112778 144764
rect 130378 144752 130384 144764
rect 112772 144724 130384 144752
rect 112772 144712 112778 144724
rect 130378 144712 130384 144724
rect 130436 144712 130442 144764
rect 173802 144712 173808 144764
rect 173860 144752 173866 144764
rect 194962 144752 194968 144764
rect 173860 144724 194968 144752
rect 173860 144712 173866 144724
rect 194962 144712 194968 144724
rect 195020 144712 195026 144764
rect 110782 144644 110788 144696
rect 110840 144684 110846 144696
rect 130562 144684 130568 144696
rect 110840 144656 130568 144684
rect 110840 144644 110846 144656
rect 130562 144644 130568 144656
rect 130620 144644 130626 144696
rect 169662 144644 169668 144696
rect 169720 144684 169726 144696
rect 196250 144684 196256 144696
rect 169720 144656 196256 144684
rect 169720 144644 169726 144656
rect 196250 144644 196256 144656
rect 196308 144644 196314 144696
rect 114002 144576 114008 144628
rect 114060 144616 114066 144628
rect 137002 144616 137008 144628
rect 114060 144588 137008 144616
rect 114060 144576 114066 144588
rect 137002 144576 137008 144588
rect 137060 144576 137066 144628
rect 165522 144576 165528 144628
rect 165580 144616 165586 144628
rect 193582 144616 193588 144628
rect 165580 144588 193588 144616
rect 165580 144576 165586 144588
rect 193582 144576 193588 144588
rect 193640 144576 193646 144628
rect 116486 144508 116492 144560
rect 116544 144548 116550 144560
rect 144178 144548 144184 144560
rect 116544 144520 144184 144548
rect 116544 144508 116550 144520
rect 144178 144508 144184 144520
rect 144236 144508 144242 144560
rect 160094 144508 160100 144560
rect 160152 144548 160158 144560
rect 194226 144548 194232 144560
rect 160152 144520 194232 144548
rect 160152 144508 160158 144520
rect 194226 144508 194232 144520
rect 194284 144508 194290 144560
rect 113910 144440 113916 144492
rect 113968 144480 113974 144492
rect 142522 144480 142528 144492
rect 113968 144452 142528 144480
rect 113968 144440 113974 144452
rect 142522 144440 142528 144452
rect 142580 144440 142586 144492
rect 162486 144440 162492 144492
rect 162544 144480 162550 144492
rect 193398 144480 193404 144492
rect 162544 144452 193404 144480
rect 162544 144440 162550 144452
rect 193398 144440 193404 144452
rect 193456 144440 193462 144492
rect 119706 144372 119712 144424
rect 119764 144412 119770 144424
rect 152458 144412 152464 144424
rect 119764 144384 152464 144412
rect 119764 144372 119770 144384
rect 152458 144372 152464 144384
rect 152516 144372 152522 144424
rect 159450 144372 159456 144424
rect 159508 144412 159514 144424
rect 193674 144412 193680 144424
rect 159508 144384 193680 144412
rect 159508 144372 159514 144384
rect 193674 144372 193680 144384
rect 193732 144372 193738 144424
rect 117866 144304 117872 144356
rect 117924 144344 117930 144356
rect 151906 144344 151912 144356
rect 117924 144316 151912 144344
rect 117924 144304 117930 144316
rect 151906 144304 151912 144316
rect 151964 144304 151970 144356
rect 154482 144304 154488 144356
rect 154540 144344 154546 144356
rect 188246 144344 188252 144356
rect 154540 144316 188252 144344
rect 154540 144304 154546 144316
rect 188246 144304 188252 144316
rect 188304 144304 188310 144356
rect 111058 144236 111064 144288
rect 111116 144276 111122 144288
rect 131206 144276 131212 144288
rect 111116 144248 131212 144276
rect 111116 144236 111122 144248
rect 131206 144236 131212 144248
rect 131264 144276 131270 144288
rect 188522 144276 188528 144288
rect 131264 144248 188528 144276
rect 131264 144236 131270 144248
rect 188522 144236 188528 144248
rect 188580 144236 188586 144288
rect 118234 144168 118240 144220
rect 118292 144208 118298 144220
rect 130194 144208 130200 144220
rect 118292 144180 130200 144208
rect 118292 144168 118298 144180
rect 130194 144168 130200 144180
rect 130252 144208 130258 144220
rect 189718 144208 189724 144220
rect 130252 144180 189724 144208
rect 130252 144168 130258 144180
rect 189718 144168 189724 144180
rect 189776 144168 189782 144220
rect 180334 144100 180340 144152
rect 180392 144140 180398 144152
rect 191282 144140 191288 144152
rect 180392 144112 191288 144140
rect 180392 144100 180398 144112
rect 191282 144100 191288 144112
rect 191340 144100 191346 144152
rect 118326 143556 118332 143608
rect 118384 143596 118390 143608
rect 145282 143596 145288 143608
rect 118384 143568 145288 143596
rect 118384 143556 118390 143568
rect 145282 143556 145288 143568
rect 145340 143556 145346 143608
rect 116670 143488 116676 143540
rect 116728 143528 116734 143540
rect 128446 143528 128452 143540
rect 116728 143500 128452 143528
rect 116728 143488 116734 143500
rect 128446 143488 128452 143500
rect 128504 143488 128510 143540
rect 128906 143488 128912 143540
rect 128964 143528 128970 143540
rect 580350 143528 580356 143540
rect 128964 143500 580356 143528
rect 128964 143488 128970 143500
rect 580350 143488 580356 143500
rect 580408 143488 580414 143540
rect 114002 143420 114008 143472
rect 114060 143460 114066 143472
rect 127710 143460 127716 143472
rect 114060 143432 127716 143460
rect 114060 143420 114066 143432
rect 127710 143420 127716 143432
rect 127768 143420 127774 143472
rect 129734 143420 129740 143472
rect 129792 143460 129798 143472
rect 137554 143460 137560 143472
rect 129792 143432 137560 143460
rect 129792 143420 129798 143432
rect 137554 143420 137560 143432
rect 137612 143420 137618 143472
rect 146294 143420 146300 143472
rect 146352 143460 146358 143472
rect 149146 143460 149152 143472
rect 146352 143432 149152 143460
rect 146352 143420 146358 143432
rect 149146 143420 149152 143432
rect 149204 143420 149210 143472
rect 176286 143420 176292 143472
rect 176344 143460 176350 143472
rect 179138 143460 179144 143472
rect 176344 143432 179144 143460
rect 176344 143420 176350 143432
rect 179138 143420 179144 143432
rect 179196 143420 179202 143472
rect 180426 143420 180432 143472
rect 180484 143460 180490 143472
rect 191466 143460 191472 143472
rect 180484 143432 191472 143460
rect 180484 143420 180490 143432
rect 191466 143420 191472 143432
rect 191524 143420 191530 143472
rect 118418 143352 118424 143404
rect 118476 143392 118482 143404
rect 133138 143392 133144 143404
rect 118476 143364 133144 143392
rect 118476 143352 118482 143364
rect 133138 143352 133144 143364
rect 133196 143352 133202 143404
rect 172882 143352 172888 143404
rect 172940 143392 172946 143404
rect 179322 143392 179328 143404
rect 172940 143364 179328 143392
rect 172940 143352 172946 143364
rect 179322 143352 179328 143364
rect 179380 143352 179386 143404
rect 185670 143352 185676 143404
rect 185728 143392 185734 143404
rect 196618 143392 196624 143404
rect 185728 143364 196624 143392
rect 185728 143352 185734 143364
rect 196618 143352 196624 143364
rect 196676 143352 196682 143404
rect 116578 143284 116584 143336
rect 116636 143324 116642 143336
rect 131482 143324 131488 143336
rect 116636 143296 131488 143324
rect 116636 143284 116642 143296
rect 131482 143284 131488 143296
rect 131540 143284 131546 143336
rect 131574 143284 131580 143336
rect 131632 143324 131638 143336
rect 135438 143324 135444 143336
rect 131632 143296 135444 143324
rect 131632 143284 131638 143296
rect 135438 143284 135444 143296
rect 135496 143284 135502 143336
rect 171042 143284 171048 143336
rect 171100 143324 171106 143336
rect 178402 143324 178408 143336
rect 171100 143296 178408 143324
rect 171100 143284 171106 143296
rect 178402 143284 178408 143296
rect 178460 143284 178466 143336
rect 181530 143284 181536 143336
rect 181588 143324 181594 143336
rect 190086 143324 190092 143336
rect 181588 143296 190092 143324
rect 181588 143284 181594 143296
rect 190086 143284 190092 143296
rect 190144 143284 190150 143336
rect 190178 143284 190184 143336
rect 190236 143324 190242 143336
rect 198366 143324 198372 143336
rect 190236 143296 198372 143324
rect 190236 143284 190242 143296
rect 198366 143284 198372 143296
rect 198424 143284 198430 143336
rect 116762 143216 116768 143268
rect 116820 143256 116826 143268
rect 134794 143256 134800 143268
rect 116820 143228 134800 143256
rect 116820 143216 116826 143228
rect 134794 143216 134800 143228
rect 134852 143216 134858 143268
rect 175734 143216 175740 143268
rect 175792 143256 175798 143268
rect 179414 143256 179420 143268
rect 175792 143228 179420 143256
rect 175792 143216 175798 143228
rect 179414 143216 179420 143228
rect 179472 143216 179478 143268
rect 183738 143216 183744 143268
rect 183796 143256 183802 143268
rect 197814 143256 197820 143268
rect 183796 143228 197820 143256
rect 183796 143216 183802 143228
rect 197814 143216 197820 143228
rect 197872 143216 197878 143268
rect 118142 143148 118148 143200
rect 118200 143188 118206 143200
rect 136634 143188 136640 143200
rect 118200 143160 136640 143188
rect 118200 143148 118206 143160
rect 136634 143148 136640 143160
rect 136692 143148 136698 143200
rect 176562 143148 176568 143200
rect 176620 143188 176626 143200
rect 192386 143188 192392 143200
rect 176620 143160 192392 143188
rect 176620 143148 176626 143160
rect 192386 143148 192392 143160
rect 192444 143148 192450 143200
rect 120902 143080 120908 143132
rect 120960 143120 120966 143132
rect 141602 143120 141608 143132
rect 120960 143092 141608 143120
rect 120960 143080 120966 143092
rect 141602 143080 141608 143092
rect 141660 143080 141666 143132
rect 170214 143080 170220 143132
rect 170272 143120 170278 143132
rect 191190 143120 191196 143132
rect 170272 143092 191196 143120
rect 170272 143080 170278 143092
rect 191190 143080 191196 143092
rect 191248 143080 191254 143132
rect 119522 143012 119528 143064
rect 119580 143052 119586 143064
rect 139762 143052 139768 143064
rect 119580 143024 139768 143052
rect 119580 143012 119586 143024
rect 139762 143012 139768 143024
rect 139820 143012 139826 143064
rect 168282 143012 168288 143064
rect 168340 143052 168346 143064
rect 184106 143052 184112 143064
rect 168340 143024 184112 143052
rect 168340 143012 168346 143024
rect 184106 143012 184112 143024
rect 184164 143012 184170 143064
rect 184290 143012 184296 143064
rect 184348 143052 184354 143064
rect 190178 143052 190184 143064
rect 184348 143024 190184 143052
rect 184348 143012 184354 143024
rect 190178 143012 190184 143024
rect 190236 143012 190242 143064
rect 119614 142944 119620 142996
rect 119672 142984 119678 142996
rect 143074 142984 143080 142996
rect 119672 142956 143080 142984
rect 119672 142944 119678 142956
rect 143074 142944 143080 142956
rect 143132 142944 143138 142996
rect 174630 142944 174636 142996
rect 174688 142984 174694 142996
rect 197630 142984 197636 142996
rect 174688 142956 197636 142984
rect 174688 142944 174694 142956
rect 197630 142944 197636 142956
rect 197688 142944 197694 142996
rect 111242 142876 111248 142928
rect 111300 142916 111306 142928
rect 134242 142916 134248 142928
rect 111300 142888 134248 142916
rect 111300 142876 111306 142888
rect 134242 142876 134248 142888
rect 134300 142876 134306 142928
rect 166902 142876 166908 142928
rect 166960 142916 166966 142928
rect 191006 142916 191012 142928
rect 166960 142888 191012 142916
rect 166960 142876 166966 142888
rect 191006 142876 191012 142888
rect 191064 142876 191070 142928
rect 108114 142808 108120 142860
rect 108172 142848 108178 142860
rect 116486 142848 116492 142860
rect 108172 142820 116492 142848
rect 108172 142808 108178 142820
rect 116486 142808 116492 142820
rect 116544 142808 116550 142860
rect 120994 142808 121000 142860
rect 121052 142848 121058 142860
rect 151354 142848 151360 142860
rect 121052 142820 151360 142848
rect 121052 142808 121058 142820
rect 151354 142808 151360 142820
rect 151412 142808 151418 142860
rect 158622 142808 158628 142860
rect 158680 142848 158686 142860
rect 191098 142848 191104 142860
rect 158680 142820 191104 142848
rect 158680 142808 158686 142820
rect 191098 142808 191104 142820
rect 191156 142808 191162 142860
rect 118326 142740 118332 142792
rect 118384 142780 118390 142792
rect 118384 142752 126652 142780
rect 118384 142740 118390 142752
rect 112622 142672 112628 142724
rect 112680 142712 112686 142724
rect 124306 142712 124312 142724
rect 112680 142684 124312 142712
rect 112680 142672 112686 142684
rect 124306 142672 124312 142684
rect 124364 142672 124370 142724
rect 126624 142712 126652 142752
rect 129826 142740 129832 142792
rect 129884 142780 129890 142792
rect 135898 142780 135904 142792
rect 129884 142752 135904 142780
rect 129884 142740 129890 142752
rect 135898 142740 135904 142752
rect 135956 142740 135962 142792
rect 178126 142740 178132 142792
rect 178184 142780 178190 142792
rect 178586 142780 178592 142792
rect 178184 142752 178592 142780
rect 178184 142740 178190 142752
rect 178586 142740 178592 142752
rect 178644 142740 178650 142792
rect 184106 142740 184112 142792
rect 184164 142780 184170 142792
rect 189626 142780 189632 142792
rect 184164 142752 189632 142780
rect 184164 142740 184170 142752
rect 189626 142740 189632 142752
rect 189684 142740 189690 142792
rect 130470 142712 130476 142724
rect 126624 142684 130476 142712
rect 130470 142672 130476 142684
rect 130528 142672 130534 142724
rect 177390 142672 177396 142724
rect 177448 142712 177454 142724
rect 179506 142712 179512 142724
rect 177448 142684 179512 142712
rect 177448 142672 177454 142684
rect 179506 142672 179512 142684
rect 179564 142672 179570 142724
rect 178218 142536 178224 142588
rect 178276 142576 178282 142588
rect 187694 142576 187700 142588
rect 178276 142548 187700 142576
rect 178276 142536 178282 142548
rect 187694 142536 187700 142548
rect 187752 142536 187758 142588
rect 129918 142196 129924 142248
rect 129976 142236 129982 142248
rect 133874 142236 133880 142248
rect 129976 142208 133880 142236
rect 129976 142196 129982 142208
rect 133874 142196 133880 142208
rect 133932 142196 133938 142248
rect 155586 142196 155592 142248
rect 155644 142236 155650 142248
rect 157334 142236 157340 142248
rect 155644 142208 157340 142236
rect 155644 142196 155650 142208
rect 157334 142196 157340 142208
rect 157392 142196 157398 142248
rect 159174 142196 159180 142248
rect 159232 142236 159238 142248
rect 161474 142236 161480 142248
rect 159232 142208 161480 142236
rect 159232 142196 159238 142208
rect 161474 142196 161480 142208
rect 161532 142196 161538 142248
rect 3418 142128 3424 142180
rect 3476 142168 3482 142180
rect 183738 142168 183744 142180
rect 3476 142140 183744 142168
rect 3476 142128 3482 142140
rect 183738 142128 183744 142140
rect 183796 142128 183802 142180
rect 120718 142060 120724 142112
rect 120776 142100 120782 142112
rect 126054 142100 126060 142112
rect 120776 142072 126060 142100
rect 120776 142060 120782 142072
rect 126054 142060 126060 142072
rect 126112 142060 126118 142112
rect 157334 142060 157340 142112
rect 157392 142100 157398 142112
rect 189442 142100 189448 142112
rect 157392 142072 189448 142100
rect 157392 142060 157398 142072
rect 189442 142060 189448 142072
rect 189500 142060 189506 142112
rect 117958 141924 117964 141976
rect 118016 141964 118022 141976
rect 126790 141964 126796 141976
rect 118016 141936 126796 141964
rect 118016 141924 118022 141936
rect 126790 141924 126796 141936
rect 126848 141924 126854 141976
rect 184198 141924 184204 141976
rect 184256 141964 184262 141976
rect 187234 141964 187240 141976
rect 184256 141936 187240 141964
rect 184256 141924 184262 141936
rect 187234 141924 187240 141936
rect 187292 141924 187298 141976
rect 183186 141856 183192 141908
rect 183244 141896 183250 141908
rect 193766 141896 193772 141908
rect 183244 141868 193772 141896
rect 183244 141856 183250 141868
rect 193766 141856 193772 141868
rect 193824 141856 193830 141908
rect 115474 141788 115480 141840
rect 115532 141828 115538 141840
rect 127342 141828 127348 141840
rect 115532 141800 127348 141828
rect 115532 141788 115538 141800
rect 127342 141788 127348 141800
rect 127400 141788 127406 141840
rect 181990 141788 181996 141840
rect 182048 141828 182054 141840
rect 196342 141828 196348 141840
rect 182048 141800 196348 141828
rect 182048 141788 182054 141800
rect 196342 141788 196348 141800
rect 196400 141788 196406 141840
rect 114094 141720 114100 141772
rect 114152 141760 114158 141772
rect 126238 141760 126244 141772
rect 114152 141732 126244 141760
rect 114152 141720 114158 141732
rect 126238 141720 126244 141732
rect 126296 141720 126302 141772
rect 179506 141720 179512 141772
rect 179564 141760 179570 141772
rect 180334 141760 180340 141772
rect 179564 141732 180340 141760
rect 179564 141720 179570 141732
rect 180334 141720 180340 141732
rect 180392 141760 180398 141772
rect 197722 141760 197728 141772
rect 180392 141732 197728 141760
rect 180392 141720 180398 141732
rect 197722 141720 197728 141732
rect 197780 141720 197786 141772
rect 119890 141652 119896 141704
rect 119948 141692 119954 141704
rect 138106 141692 138112 141704
rect 119948 141664 138112 141692
rect 119948 141652 119954 141664
rect 138106 141652 138112 141664
rect 138164 141652 138170 141704
rect 175182 141652 175188 141704
rect 175240 141692 175246 141704
rect 193490 141692 193496 141704
rect 175240 141664 193496 141692
rect 175240 141652 175246 141664
rect 193490 141652 193496 141664
rect 193548 141652 193554 141704
rect 118142 141584 118148 141636
rect 118200 141624 118206 141636
rect 146846 141624 146852 141636
rect 118200 141596 146852 141624
rect 118200 141584 118206 141596
rect 146846 141584 146852 141596
rect 146904 141584 146910 141636
rect 170766 141584 170772 141636
rect 170824 141624 170830 141636
rect 192018 141624 192024 141636
rect 170824 141596 192024 141624
rect 170824 141584 170830 141596
rect 192018 141584 192024 141596
rect 192076 141584 192082 141636
rect 120810 141516 120816 141568
rect 120868 141556 120874 141568
rect 152366 141556 152372 141568
rect 120868 141528 152372 141556
rect 120868 141516 120874 141528
rect 152366 141516 152372 141528
rect 152424 141516 152430 141568
rect 169110 141516 169116 141568
rect 169168 141556 169174 141568
rect 192294 141556 192300 141568
rect 169168 141528 192300 141556
rect 169168 141516 169174 141528
rect 192294 141516 192300 141528
rect 192352 141516 192358 141568
rect 120902 141448 120908 141500
rect 120960 141488 120966 141500
rect 153286 141488 153292 141500
rect 120960 141460 153292 141488
rect 120960 141448 120966 141460
rect 153286 141448 153292 141460
rect 153344 141448 153350 141500
rect 167454 141448 167460 141500
rect 167512 141488 167518 141500
rect 192202 141488 192208 141500
rect 167512 141460 192208 141488
rect 167512 141448 167518 141460
rect 192202 141448 192208 141460
rect 192260 141448 192266 141500
rect 119430 141380 119436 141432
rect 119488 141420 119494 141432
rect 153746 141420 153752 141432
rect 119488 141392 153752 141420
rect 119488 141380 119494 141392
rect 153746 141380 153752 141392
rect 153804 141380 153810 141432
rect 157150 141380 157156 141432
rect 157208 141420 157214 141432
rect 189350 141420 189356 141432
rect 157208 141392 189356 141420
rect 157208 141380 157214 141392
rect 189350 141380 189356 141392
rect 189408 141380 189414 141432
rect 119798 141312 119804 141364
rect 119856 141352 119862 141364
rect 123478 141352 123484 141364
rect 119856 141324 123484 141352
rect 119856 141312 119862 141324
rect 123478 141312 123484 141324
rect 123536 141312 123542 141364
rect 116854 141244 116860 141296
rect 116912 141284 116918 141296
rect 125502 141284 125508 141296
rect 116912 141256 125508 141284
rect 116912 141244 116918 141256
rect 125502 141244 125508 141256
rect 125560 141244 125566 141296
rect 185026 141176 185032 141228
rect 185084 141216 185090 141228
rect 185670 141216 185676 141228
rect 185084 141188 185676 141216
rect 185084 141176 185090 141188
rect 185670 141176 185676 141188
rect 185728 141176 185734 141228
rect 126054 141108 126060 141160
rect 126112 141148 126118 141160
rect 129458 141148 129464 141160
rect 126112 141120 129464 141148
rect 126112 141108 126118 141120
rect 129458 141108 129464 141120
rect 129516 141108 129522 141160
rect 184750 141108 184756 141160
rect 184808 141148 184814 141160
rect 190914 141148 190920 141160
rect 184808 141120 190920 141148
rect 184808 141108 184814 141120
rect 190914 141108 190920 141120
rect 190972 141108 190978 141160
rect 117958 141040 117964 141092
rect 118016 141080 118022 141092
rect 179506 141080 179512 141092
rect 118016 141052 179512 141080
rect 118016 141040 118022 141052
rect 179506 141040 179512 141052
rect 179564 141040 179570 141092
rect 17218 140972 17224 141024
rect 17276 141012 17282 141024
rect 185026 141012 185032 141024
rect 17276 140984 185032 141012
rect 17276 140972 17282 140984
rect 185026 140972 185032 140984
rect 185084 140972 185090 141024
rect 8938 140904 8944 140956
rect 8996 140944 9002 140956
rect 182910 140944 182916 140956
rect 8996 140916 182916 140944
rect 8996 140904 9002 140916
rect 182910 140904 182916 140916
rect 182968 140904 182974 140956
rect 185854 140904 185860 140956
rect 185912 140944 185918 140956
rect 191190 140944 191196 140956
rect 185912 140916 191196 140944
rect 185912 140904 185918 140916
rect 191190 140904 191196 140916
rect 191248 140904 191254 140956
rect 126790 140836 126796 140888
rect 126848 140876 126854 140888
rect 126848 140848 129320 140876
rect 126848 140836 126854 140848
rect 129292 140808 129320 140848
rect 129458 140836 129464 140888
rect 129516 140876 129522 140888
rect 327718 140876 327724 140888
rect 129516 140848 327724 140876
rect 129516 140836 129522 140848
rect 327718 140836 327724 140848
rect 327776 140836 327782 140888
rect 464338 140808 464344 140820
rect 129292 140780 464344 140808
rect 464338 140768 464344 140780
rect 464396 140768 464402 140820
rect 119522 140700 119528 140752
rect 119580 140740 119586 140752
rect 119580 140712 124996 140740
rect 119580 140700 119586 140712
rect 119338 140632 119344 140684
rect 119396 140672 119402 140684
rect 124766 140672 124772 140684
rect 119396 140644 124772 140672
rect 119396 140632 119402 140644
rect 124766 140632 124772 140644
rect 124824 140632 124830 140684
rect 124968 140672 124996 140712
rect 128354 140700 128360 140752
rect 128412 140740 128418 140752
rect 129274 140740 129280 140752
rect 128412 140712 129280 140740
rect 128412 140700 128418 140712
rect 129274 140700 129280 140712
rect 129332 140700 129338 140752
rect 131298 140700 131304 140752
rect 131356 140740 131362 140752
rect 132310 140740 132316 140752
rect 131356 140712 132316 140740
rect 131356 140700 131362 140712
rect 132310 140700 132316 140712
rect 132368 140700 132374 140752
rect 146938 140740 146944 140752
rect 142126 140712 146944 140740
rect 128998 140672 129004 140684
rect 124968 140644 129004 140672
rect 128998 140632 129004 140644
rect 129056 140632 129062 140684
rect 113634 140564 113640 140616
rect 113692 140604 113698 140616
rect 129090 140604 129096 140616
rect 113692 140576 129096 140604
rect 113692 140564 113698 140576
rect 129090 140564 129096 140576
rect 129148 140564 129154 140616
rect 120994 140496 121000 140548
rect 121052 140536 121058 140548
rect 142126 140536 142154 140712
rect 146938 140700 146944 140712
rect 146996 140700 147002 140752
rect 178034 140700 178040 140752
rect 178092 140740 178098 140752
rect 178954 140740 178960 140752
rect 178092 140712 178960 140740
rect 178092 140700 178098 140712
rect 178954 140700 178960 140712
rect 179012 140700 179018 140752
rect 190822 140740 190828 140752
rect 180766 140712 190828 140740
rect 146754 140632 146760 140684
rect 146812 140632 146818 140684
rect 173894 140632 173900 140684
rect 173952 140672 173958 140684
rect 179138 140672 179144 140684
rect 173952 140644 179144 140672
rect 173952 140632 173958 140644
rect 179138 140632 179144 140644
rect 179196 140632 179202 140684
rect 121052 140508 142154 140536
rect 121052 140496 121058 140508
rect 119246 140428 119252 140480
rect 119304 140468 119310 140480
rect 146772 140468 146800 140632
rect 171134 140564 171140 140616
rect 171192 140604 171198 140616
rect 180766 140604 180794 140712
rect 190822 140700 190828 140712
rect 190880 140700 190886 140752
rect 171192 140576 180794 140604
rect 171192 140564 171198 140576
rect 184474 140564 184480 140616
rect 184532 140604 184538 140616
rect 193950 140604 193956 140616
rect 184532 140576 193956 140604
rect 184532 140564 184538 140576
rect 193950 140564 193956 140576
rect 194008 140564 194014 140616
rect 178126 140496 178132 140548
rect 178184 140536 178190 140548
rect 178586 140536 178592 140548
rect 178184 140508 178592 140536
rect 178184 140496 178190 140508
rect 178586 140496 178592 140508
rect 178644 140496 178650 140548
rect 179966 140496 179972 140548
rect 180024 140536 180030 140548
rect 193582 140536 193588 140548
rect 180024 140508 193588 140536
rect 180024 140496 180030 140508
rect 193582 140496 193588 140508
rect 193640 140496 193646 140548
rect 119304 140440 146800 140468
rect 119304 140428 119310 140440
rect 179046 140428 179052 140480
rect 179104 140468 179110 140480
rect 196618 140468 196624 140480
rect 179104 140440 196624 140468
rect 179104 140428 179110 140440
rect 196618 140428 196624 140440
rect 196676 140428 196682 140480
rect 119430 140360 119436 140412
rect 119488 140400 119494 140412
rect 148226 140400 148232 140412
rect 119488 140372 148232 140400
rect 119488 140360 119494 140372
rect 148226 140360 148232 140372
rect 148284 140360 148290 140412
rect 171226 140360 171232 140412
rect 171284 140400 171290 140412
rect 189718 140400 189724 140412
rect 171284 140372 189724 140400
rect 171284 140360 171290 140372
rect 189718 140360 189724 140372
rect 189776 140360 189782 140412
rect 116394 140292 116400 140344
rect 116452 140332 116458 140344
rect 145558 140332 145564 140344
rect 116452 140304 145564 140332
rect 116452 140292 116458 140304
rect 145558 140292 145564 140304
rect 145616 140292 145622 140344
rect 169846 140292 169852 140344
rect 169904 140332 169910 140344
rect 189534 140332 189540 140344
rect 169904 140304 189540 140332
rect 169904 140292 169910 140304
rect 189534 140292 189540 140304
rect 189592 140292 189598 140344
rect 116578 140224 116584 140276
rect 116636 140264 116642 140276
rect 147950 140264 147956 140276
rect 116636 140236 147956 140264
rect 116636 140224 116642 140236
rect 147950 140224 147956 140236
rect 148008 140224 148014 140276
rect 171318 140224 171324 140276
rect 171376 140264 171382 140276
rect 192386 140264 192392 140276
rect 171376 140236 192392 140264
rect 171376 140224 171382 140236
rect 192386 140224 192392 140236
rect 192444 140224 192450 140276
rect 117866 140156 117872 140208
rect 117924 140196 117930 140208
rect 149422 140196 149428 140208
rect 117924 140168 149428 140196
rect 117924 140156 117930 140168
rect 149422 140156 149428 140168
rect 149480 140156 149486 140208
rect 169938 140156 169944 140208
rect 169996 140196 170002 140208
rect 185578 140196 185584 140208
rect 169996 140168 185584 140196
rect 169996 140156 170002 140168
rect 185578 140156 185584 140168
rect 185636 140156 185642 140208
rect 192570 140196 192576 140208
rect 190426 140168 192576 140196
rect 116762 140088 116768 140140
rect 116820 140128 116826 140140
rect 150066 140128 150072 140140
rect 116820 140100 150072 140128
rect 116820 140088 116826 140100
rect 150066 140088 150072 140100
rect 150124 140088 150130 140140
rect 170858 140088 170864 140140
rect 170916 140128 170922 140140
rect 190426 140128 190454 140168
rect 192570 140156 192576 140168
rect 192628 140156 192634 140208
rect 170916 140100 190454 140128
rect 170916 140088 170922 140100
rect 119154 140020 119160 140072
rect 119212 140060 119218 140072
rect 126146 140060 126152 140072
rect 119212 140032 126152 140060
rect 119212 140020 119218 140032
rect 126146 140020 126152 140032
rect 126204 140020 126210 140072
rect 126606 140020 126612 140072
rect 126664 140060 126670 140072
rect 184658 140060 184664 140072
rect 126664 140032 184664 140060
rect 126664 140020 126670 140032
rect 184658 140020 184664 140032
rect 184716 140020 184722 140072
rect 185670 140020 185676 140072
rect 185728 140060 185734 140072
rect 196434 140060 196440 140072
rect 185728 140032 196440 140060
rect 185728 140020 185734 140032
rect 196434 140020 196440 140032
rect 196492 140020 196498 140072
rect 120626 139952 120632 140004
rect 120684 139992 120690 140004
rect 129182 139992 129188 140004
rect 120684 139964 129188 139992
rect 120684 139952 120690 139964
rect 129182 139952 129188 139964
rect 129240 139952 129246 140004
rect 129458 139952 129464 140004
rect 129516 139952 129522 140004
rect 183002 139952 183008 140004
rect 183060 139992 183066 140004
rect 189902 139992 189908 140004
rect 183060 139964 189908 139992
rect 183060 139952 183066 139964
rect 189902 139952 189908 139964
rect 189960 139952 189966 140004
rect 124766 139884 124772 139936
rect 124824 139924 124830 139936
rect 129476 139924 129504 139952
rect 124824 139896 129504 139924
rect 124824 139884 124830 139896
rect 184566 139884 184572 139936
rect 184624 139924 184630 139936
rect 189626 139924 189632 139936
rect 184624 139896 189632 139924
rect 184624 139884 184630 139896
rect 189626 139884 189632 139896
rect 189684 139884 189690 139936
rect 119798 139816 119804 139868
rect 119856 139856 119862 139868
rect 126514 139856 126520 139868
rect 119856 139828 126520 139856
rect 119856 139816 119862 139828
rect 126514 139816 126520 139828
rect 126572 139816 126578 139868
rect 185578 139816 185584 139868
rect 185636 139856 185642 139868
rect 192662 139856 192668 139868
rect 185636 139828 192668 139856
rect 185636 139816 185642 139828
rect 192662 139816 192668 139828
rect 192720 139816 192726 139868
rect 118050 139680 118056 139732
rect 118108 139720 118114 139732
rect 124858 139720 124864 139732
rect 118108 139692 124864 139720
rect 118108 139680 118114 139692
rect 124858 139680 124864 139692
rect 124916 139680 124922 139732
rect 128814 139544 128820 139596
rect 128872 139584 128878 139596
rect 178034 139584 178040 139596
rect 128872 139556 178040 139584
rect 128872 139544 128878 139556
rect 178034 139544 178040 139556
rect 178092 139544 178098 139596
rect 181622 139544 181628 139596
rect 181680 139584 181686 139596
rect 188614 139584 188620 139596
rect 181680 139556 188620 139584
rect 181680 139544 181686 139556
rect 188614 139544 188620 139556
rect 188672 139544 188678 139596
rect 127526 139476 127532 139528
rect 127584 139516 127590 139528
rect 181806 139516 181812 139528
rect 127584 139488 181812 139516
rect 127584 139476 127590 139488
rect 181806 139476 181812 139488
rect 181864 139476 181870 139528
rect 124858 139408 124864 139460
rect 124916 139448 124922 139460
rect 181898 139448 181904 139460
rect 124916 139420 181904 139448
rect 124916 139408 124922 139420
rect 181898 139408 181904 139420
rect 181956 139408 181962 139460
rect 183278 139408 183284 139460
rect 183336 139448 183342 139460
rect 189810 139448 189816 139460
rect 183336 139420 189816 139448
rect 183336 139408 183342 139420
rect 189810 139408 189816 139420
rect 189868 139408 189874 139460
rect 126146 139340 126152 139392
rect 126204 139380 126210 139392
rect 126422 139380 126428 139392
rect 126204 139352 126428 139380
rect 126204 139340 126210 139352
rect 126422 139340 126428 139352
rect 126480 139340 126486 139392
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 117958 137952 117964 137964
rect 3568 137924 117964 137952
rect 3568 137912 3574 137924
rect 117958 137912 117964 137924
rect 118016 137912 118022 137964
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 31018 111772 31024 111784
rect 3200 111744 31024 111772
rect 3200 111732 3206 111744
rect 31018 111732 31024 111744
rect 31076 111732 31082 111784
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 120534 97968 120540 97980
rect 3568 97940 120540 97968
rect 3568 97928 3574 97940
rect 120534 97928 120540 97940
rect 120592 97928 120598 97980
rect 107286 89088 107292 89140
rect 107344 89088 107350 89140
rect 107304 88924 107332 89088
rect 107378 88924 107384 88936
rect 107304 88896 107384 88924
rect 107378 88884 107384 88896
rect 107436 88884 107442 88936
rect 464338 86912 464344 86964
rect 464396 86952 464402 86964
rect 580166 86952 580172 86964
rect 464396 86924 580172 86952
rect 464396 86912 464402 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 121914 81200 121920 81252
rect 121972 81240 121978 81252
rect 122190 81240 122196 81252
rect 121972 81212 122196 81240
rect 121972 81200 121978 81212
rect 122190 81200 122196 81212
rect 122248 81200 122254 81252
rect 187418 81240 187424 81252
rect 158686 81212 187424 81240
rect 124186 81144 131896 81172
rect 123110 81064 123116 81116
rect 123168 81104 123174 81116
rect 124186 81104 124214 81144
rect 123168 81076 124214 81104
rect 123168 81064 123174 81076
rect 121638 80996 121644 81048
rect 121696 81036 121702 81048
rect 121696 81008 124214 81036
rect 121696 80996 121702 81008
rect 108298 80860 108304 80912
rect 108356 80900 108362 80912
rect 120718 80900 120724 80912
rect 108356 80872 120724 80900
rect 108356 80860 108362 80872
rect 120718 80860 120724 80872
rect 120776 80860 120782 80912
rect 124186 80832 124214 81008
rect 115906 80804 123616 80832
rect 124186 80804 131804 80832
rect 115906 80764 115934 80804
rect 113146 80736 115934 80764
rect 123588 80764 123616 80804
rect 123588 80736 131712 80764
rect 71774 80656 71780 80708
rect 71832 80696 71838 80708
rect 108390 80696 108396 80708
rect 71832 80668 108396 80696
rect 71832 80656 71838 80668
rect 108390 80656 108396 80668
rect 108448 80696 108454 80708
rect 113146 80696 113174 80736
rect 131684 80708 131712 80736
rect 108448 80668 113174 80696
rect 108448 80656 108454 80668
rect 116578 80656 116584 80708
rect 116636 80696 116642 80708
rect 116636 80668 118694 80696
rect 116636 80656 116642 80668
rect 118666 80560 118694 80668
rect 120718 80656 120724 80708
rect 120776 80696 120782 80708
rect 130010 80696 130016 80708
rect 120776 80668 130016 80696
rect 120776 80656 120782 80668
rect 130010 80656 130016 80668
rect 130068 80656 130074 80708
rect 131666 80656 131672 80708
rect 131724 80656 131730 80708
rect 131776 80628 131804 80804
rect 131868 80708 131896 81144
rect 158686 81104 158714 81212
rect 187418 81200 187424 81212
rect 187476 81200 187482 81252
rect 154546 81076 158714 81104
rect 154546 80968 154574 81076
rect 187510 81064 187516 81116
rect 187568 81104 187574 81116
rect 192662 81104 192668 81116
rect 187568 81076 192668 81104
rect 187568 81064 187574 81076
rect 192662 81064 192668 81076
rect 192720 81064 192726 81116
rect 186774 81036 186780 81048
rect 151786 80940 154574 80968
rect 158686 81008 159174 81036
rect 131850 80656 131856 80708
rect 131908 80656 131914 80708
rect 132328 80668 146294 80696
rect 132328 80628 132356 80668
rect 131776 80600 132356 80628
rect 146266 80628 146294 80668
rect 146266 80600 149238 80628
rect 118666 80532 124214 80560
rect 124186 80492 124214 80532
rect 146266 80532 148870 80560
rect 146266 80492 146294 80532
rect 124186 80464 146294 80492
rect 106734 80384 106740 80436
rect 106792 80424 106798 80436
rect 107010 80424 107016 80436
rect 106792 80396 107016 80424
rect 106792 80384 106798 80396
rect 107010 80384 107016 80396
rect 107068 80384 107074 80436
rect 130746 80316 130752 80368
rect 130804 80356 130810 80368
rect 130804 80328 145006 80356
rect 130804 80316 130810 80328
rect 107010 80248 107016 80300
rect 107068 80288 107074 80300
rect 107194 80288 107200 80300
rect 107068 80260 107200 80288
rect 107068 80248 107074 80260
rect 107194 80248 107200 80260
rect 107252 80248 107258 80300
rect 131850 80248 131856 80300
rect 131908 80288 131914 80300
rect 131908 80260 143626 80288
rect 131908 80248 131914 80260
rect 131758 80180 131764 80232
rect 131816 80220 131822 80232
rect 131816 80192 142154 80220
rect 131816 80180 131822 80192
rect 131574 80112 131580 80164
rect 131632 80152 131638 80164
rect 131632 80124 134978 80152
rect 131632 80112 131638 80124
rect 119154 80044 119160 80096
rect 119212 80084 119218 80096
rect 130746 80084 130752 80096
rect 119212 80056 130752 80084
rect 119212 80044 119218 80056
rect 130746 80044 130752 80056
rect 130804 80044 130810 80096
rect 131666 80044 131672 80096
rect 131724 80084 131730 80096
rect 131724 80056 134886 80084
rect 131724 80044 131730 80056
rect 130654 79976 130660 80028
rect 130712 80016 130718 80028
rect 130712 79988 133322 80016
rect 130712 79976 130718 79988
rect 133294 79960 133322 79988
rect 130470 79908 130476 79960
rect 130528 79948 130534 79960
rect 132632 79948 132638 79960
rect 130528 79920 132638 79948
rect 130528 79908 130534 79920
rect 132632 79908 132638 79920
rect 132690 79908 132696 79960
rect 132816 79908 132822 79960
rect 132874 79908 132880 79960
rect 133092 79908 133098 79960
rect 133150 79908 133156 79960
rect 133276 79908 133282 79960
rect 133334 79908 133340 79960
rect 133368 79908 133374 79960
rect 133426 79908 133432 79960
rect 133460 79908 133466 79960
rect 133518 79908 133524 79960
rect 133552 79908 133558 79960
rect 133610 79948 133616 79960
rect 133610 79908 133644 79948
rect 133736 79908 133742 79960
rect 133794 79908 133800 79960
rect 133828 79908 133834 79960
rect 133886 79908 133892 79960
rect 133920 79908 133926 79960
rect 133978 79908 133984 79960
rect 134104 79908 134110 79960
rect 134162 79908 134168 79960
rect 134380 79908 134386 79960
rect 134438 79948 134444 79960
rect 134438 79908 134472 79948
rect 134564 79908 134570 79960
rect 134622 79908 134628 79960
rect 132126 79840 132132 79892
rect 132184 79880 132190 79892
rect 132834 79880 132862 79908
rect 132184 79852 132862 79880
rect 132184 79840 132190 79852
rect 132908 79840 132914 79892
rect 132966 79840 132972 79892
rect 129458 79772 129464 79824
rect 129516 79812 129522 79824
rect 132926 79812 132954 79840
rect 129516 79784 132954 79812
rect 129516 79772 129522 79784
rect 133110 79756 133138 79908
rect 133184 79840 133190 79892
rect 133242 79880 133248 79892
rect 133242 79840 133276 79880
rect 109862 79704 109868 79756
rect 109920 79744 109926 79756
rect 131758 79744 131764 79756
rect 109920 79716 131764 79744
rect 109920 79704 109926 79716
rect 131758 79704 131764 79716
rect 131816 79704 131822 79756
rect 133110 79716 133144 79756
rect 133138 79704 133144 79716
rect 133196 79704 133202 79756
rect 116210 79636 116216 79688
rect 116268 79676 116274 79688
rect 133248 79676 133276 79840
rect 133386 79756 133414 79908
rect 133478 79824 133506 79908
rect 133478 79784 133512 79824
rect 133506 79772 133512 79784
rect 133564 79772 133570 79824
rect 133386 79716 133420 79756
rect 133414 79704 133420 79716
rect 133472 79704 133478 79756
rect 133322 79676 133328 79688
rect 116268 79648 128354 79676
rect 133248 79648 133328 79676
rect 116268 79636 116274 79648
rect 112346 79568 112352 79620
rect 112404 79608 112410 79620
rect 122834 79608 122840 79620
rect 112404 79580 122840 79608
rect 112404 79568 112410 79580
rect 122834 79568 122840 79580
rect 122892 79608 122898 79620
rect 124122 79608 124128 79620
rect 122892 79580 124128 79608
rect 122892 79568 122898 79580
rect 124122 79568 124128 79580
rect 124180 79568 124186 79620
rect 113818 79500 113824 79552
rect 113876 79540 113882 79552
rect 125594 79540 125600 79552
rect 113876 79512 125600 79540
rect 113876 79500 113882 79512
rect 125594 79500 125600 79512
rect 125652 79500 125658 79552
rect 106826 79432 106832 79484
rect 106884 79472 106890 79484
rect 126238 79472 126244 79484
rect 106884 79444 126244 79472
rect 106884 79432 106890 79444
rect 126238 79432 126244 79444
rect 126296 79432 126302 79484
rect 128326 79472 128354 79648
rect 133322 79636 133328 79648
rect 133380 79636 133386 79688
rect 133046 79568 133052 79620
rect 133104 79608 133110 79620
rect 133616 79608 133644 79908
rect 133754 79824 133782 79908
rect 133736 79772 133742 79824
rect 133794 79772 133800 79824
rect 133846 79688 133874 79908
rect 133782 79636 133788 79688
rect 133840 79648 133874 79688
rect 133840 79636 133846 79648
rect 133104 79580 133644 79608
rect 133104 79568 133110 79580
rect 132402 79500 132408 79552
rect 132460 79540 132466 79552
rect 133938 79540 133966 79908
rect 134012 79840 134018 79892
rect 134070 79840 134076 79892
rect 134030 79620 134058 79840
rect 134122 79688 134150 79908
rect 134196 79840 134202 79892
rect 134254 79840 134260 79892
rect 134288 79840 134294 79892
rect 134346 79880 134352 79892
rect 134346 79840 134380 79880
rect 134214 79756 134242 79840
rect 134214 79716 134248 79756
rect 134242 79704 134248 79716
rect 134300 79704 134306 79756
rect 134122 79648 134156 79688
rect 134150 79636 134156 79648
rect 134208 79636 134214 79688
rect 134352 79676 134380 79840
rect 134444 79688 134472 79908
rect 134260 79648 134380 79676
rect 134030 79580 134064 79620
rect 134058 79568 134064 79580
rect 134116 79568 134122 79620
rect 132460 79512 133966 79540
rect 134260 79540 134288 79648
rect 134426 79636 134432 79688
rect 134484 79636 134490 79688
rect 134334 79568 134340 79620
rect 134392 79608 134398 79620
rect 134582 79608 134610 79908
rect 134748 79840 134754 79892
rect 134806 79840 134812 79892
rect 134858 79880 134886 80056
rect 134950 79960 134978 80124
rect 142126 80084 142154 80192
rect 139918 80056 141694 80084
rect 142126 80056 142706 80084
rect 135134 79988 138014 80016
rect 134932 79908 134938 79960
rect 134990 79908 134996 79960
rect 135134 79880 135162 79988
rect 137986 79960 138014 79988
rect 135208 79908 135214 79960
rect 135266 79908 135272 79960
rect 135300 79908 135306 79960
rect 135358 79908 135364 79960
rect 136128 79908 136134 79960
rect 136186 79908 136192 79960
rect 136312 79908 136318 79960
rect 136370 79948 136376 79960
rect 136370 79920 136496 79948
rect 136370 79908 136376 79920
rect 134858 79852 135162 79880
rect 134766 79620 134794 79840
rect 135226 79688 135254 79908
rect 135318 79824 135346 79908
rect 135944 79840 135950 79892
rect 136002 79880 136008 79892
rect 136002 79840 136036 79880
rect 135318 79784 135352 79824
rect 135346 79772 135352 79784
rect 135404 79772 135410 79824
rect 135668 79772 135674 79824
rect 135726 79772 135732 79824
rect 135760 79772 135766 79824
rect 135818 79812 135824 79824
rect 135818 79772 135852 79812
rect 135162 79636 135168 79688
rect 135220 79648 135254 79688
rect 135686 79688 135714 79772
rect 135686 79648 135720 79688
rect 135220 79636 135226 79648
rect 135714 79636 135720 79648
rect 135772 79636 135778 79688
rect 134392 79580 134610 79608
rect 134392 79568 134398 79580
rect 134702 79568 134708 79620
rect 134760 79580 134794 79620
rect 134760 79568 134766 79580
rect 135622 79568 135628 79620
rect 135680 79608 135686 79620
rect 135824 79608 135852 79772
rect 136008 79688 136036 79840
rect 136146 79688 136174 79908
rect 136220 79840 136226 79892
rect 136278 79880 136284 79892
rect 136278 79840 136312 79880
rect 136284 79756 136312 79840
rect 136358 79772 136364 79824
rect 136416 79772 136422 79824
rect 136266 79704 136272 79756
rect 136324 79704 136330 79756
rect 135990 79636 135996 79688
rect 136048 79636 136054 79688
rect 136146 79648 136180 79688
rect 136174 79636 136180 79648
rect 136232 79636 136238 79688
rect 135680 79580 135852 79608
rect 135680 79568 135686 79580
rect 134518 79540 134524 79552
rect 134260 79512 134524 79540
rect 132460 79500 132466 79512
rect 134518 79500 134524 79512
rect 134576 79540 134582 79552
rect 135070 79540 135076 79552
rect 134576 79512 135076 79540
rect 134576 79500 134582 79512
rect 135070 79500 135076 79512
rect 135128 79500 135134 79552
rect 135806 79500 135812 79552
rect 135864 79540 135870 79552
rect 136376 79540 136404 79772
rect 136468 79552 136496 79920
rect 136680 79908 136686 79960
rect 136738 79908 136744 79960
rect 137140 79948 137146 79960
rect 136928 79920 137146 79948
rect 136698 79756 136726 79908
rect 136698 79716 136732 79756
rect 136726 79704 136732 79716
rect 136784 79704 136790 79756
rect 136928 79744 136956 79920
rect 137140 79908 137146 79920
rect 137198 79908 137204 79960
rect 137416 79948 137422 79960
rect 137296 79920 137422 79948
rect 137094 79744 137100 79756
rect 136928 79716 137100 79744
rect 136928 79620 136956 79716
rect 137094 79704 137100 79716
rect 137152 79704 137158 79756
rect 137296 79688 137324 79920
rect 137416 79908 137422 79920
rect 137474 79908 137480 79960
rect 137968 79908 137974 79960
rect 138026 79908 138032 79960
rect 138060 79908 138066 79960
rect 138118 79908 138124 79960
rect 138152 79908 138158 79960
rect 138210 79908 138216 79960
rect 138244 79908 138250 79960
rect 138302 79908 138308 79960
rect 138612 79948 138618 79960
rect 138354 79920 138618 79948
rect 137692 79840 137698 79892
rect 137750 79840 137756 79892
rect 138078 79880 138106 79908
rect 138032 79852 138106 79880
rect 137278 79636 137284 79688
rect 137336 79636 137342 79688
rect 137554 79636 137560 79688
rect 137612 79676 137618 79688
rect 137710 79676 137738 79840
rect 138032 79824 138060 79852
rect 138170 79824 138198 79908
rect 137876 79772 137882 79824
rect 137934 79772 137940 79824
rect 138014 79772 138020 79824
rect 138072 79772 138078 79824
rect 138106 79772 138112 79824
rect 138164 79784 138198 79824
rect 138164 79772 138170 79784
rect 137894 79688 137922 79772
rect 138262 79756 138290 79908
rect 138198 79704 138204 79756
rect 138256 79716 138290 79756
rect 138256 79704 138262 79716
rect 137612 79648 137738 79676
rect 137612 79636 137618 79648
rect 137830 79636 137836 79688
rect 137888 79648 137922 79688
rect 137888 79636 137894 79648
rect 136910 79568 136916 79620
rect 136968 79568 136974 79620
rect 135864 79512 136404 79540
rect 135864 79500 135870 79512
rect 136450 79500 136456 79552
rect 136508 79500 136514 79552
rect 138354 79540 138382 79920
rect 138612 79908 138618 79920
rect 138670 79908 138676 79960
rect 139256 79948 139262 79960
rect 139228 79908 139262 79948
rect 139314 79908 139320 79960
rect 139624 79908 139630 79960
rect 139682 79908 139688 79960
rect 138796 79840 138802 79892
rect 138854 79840 138860 79892
rect 139072 79840 139078 79892
rect 139130 79880 139136 79892
rect 139130 79840 139164 79880
rect 138814 79744 138842 79840
rect 138814 79716 139072 79744
rect 138566 79540 138572 79552
rect 138354 79512 138572 79540
rect 138566 79500 138572 79512
rect 138624 79500 138630 79552
rect 139044 79540 139072 79716
rect 139136 79608 139164 79840
rect 139228 79688 139256 79908
rect 139210 79636 139216 79688
rect 139268 79636 139274 79688
rect 139302 79608 139308 79620
rect 139136 79580 139308 79608
rect 139302 79568 139308 79580
rect 139360 79568 139366 79620
rect 139394 79568 139400 79620
rect 139452 79608 139458 79620
rect 139642 79608 139670 79908
rect 139918 79620 139946 80056
rect 141666 80016 141694 80056
rect 142678 80016 142706 80056
rect 139452 79580 139670 79608
rect 139452 79568 139458 79580
rect 139854 79568 139860 79620
rect 139912 79580 139946 79620
rect 140056 79988 141602 80016
rect 141666 79988 142614 80016
rect 142678 79988 143534 80016
rect 139912 79568 139918 79580
rect 140056 79552 140084 79988
rect 141574 79960 141602 79988
rect 142586 79960 142614 79988
rect 140360 79948 140366 79960
rect 140148 79920 140366 79948
rect 139210 79540 139216 79552
rect 139044 79512 139216 79540
rect 139210 79500 139216 79512
rect 139268 79500 139274 79552
rect 140038 79500 140044 79552
rect 140096 79500 140102 79552
rect 140148 79540 140176 79920
rect 140360 79908 140366 79920
rect 140418 79908 140424 79960
rect 140452 79908 140458 79960
rect 140510 79908 140516 79960
rect 140544 79908 140550 79960
rect 140602 79908 140608 79960
rect 141464 79908 141470 79960
rect 141522 79908 141528 79960
rect 141556 79908 141562 79960
rect 141614 79908 141620 79960
rect 142292 79948 142298 79960
rect 142264 79908 142298 79948
rect 142350 79908 142356 79960
rect 142568 79908 142574 79960
rect 142626 79908 142632 79960
rect 142752 79908 142758 79960
rect 142810 79908 142816 79960
rect 143396 79908 143402 79960
rect 143454 79908 143460 79960
rect 140470 79824 140498 79908
rect 140406 79772 140412 79824
rect 140464 79784 140498 79824
rect 140464 79772 140470 79784
rect 140222 79568 140228 79620
rect 140280 79608 140286 79620
rect 140562 79608 140590 79908
rect 141004 79880 141010 79892
rect 140280 79580 140590 79608
rect 140884 79852 141010 79880
rect 140280 79568 140286 79580
rect 140884 79552 140912 79852
rect 141004 79840 141010 79852
rect 141062 79840 141068 79892
rect 141482 79620 141510 79908
rect 141648 79840 141654 79892
rect 141706 79840 141712 79892
rect 141832 79840 141838 79892
rect 141890 79880 141896 79892
rect 142016 79880 142022 79892
rect 141890 79840 141924 79880
rect 141418 79568 141424 79620
rect 141476 79580 141510 79620
rect 141476 79568 141482 79580
rect 140682 79540 140688 79552
rect 140148 79512 140688 79540
rect 140682 79500 140688 79512
rect 140740 79500 140746 79552
rect 140866 79500 140872 79552
rect 140924 79500 140930 79552
rect 141234 79500 141240 79552
rect 141292 79540 141298 79552
rect 141666 79540 141694 79840
rect 141896 79688 141924 79840
rect 141988 79840 142022 79880
rect 142074 79840 142080 79892
rect 141988 79688 142016 79840
rect 142264 79688 142292 79908
rect 142770 79756 142798 79908
rect 143028 79840 143034 79892
rect 143086 79840 143092 79892
rect 142614 79704 142620 79756
rect 142672 79704 142678 79756
rect 142770 79716 142804 79756
rect 142798 79704 142804 79716
rect 142856 79704 142862 79756
rect 143046 79744 143074 79840
rect 143414 79756 143442 79908
rect 143506 79880 143534 79988
rect 143598 79948 143626 80260
rect 143874 79988 144270 80016
rect 143672 79948 143678 79960
rect 143598 79920 143678 79948
rect 143672 79908 143678 79920
rect 143730 79908 143736 79960
rect 143874 79880 143902 79988
rect 144242 79960 144270 79988
rect 144978 79960 145006 80328
rect 146680 79988 147030 80016
rect 144132 79948 144138 79960
rect 144104 79908 144138 79948
rect 144190 79908 144196 79960
rect 144224 79908 144230 79960
rect 144282 79908 144288 79960
rect 144960 79908 144966 79960
rect 145018 79908 145024 79960
rect 145328 79908 145334 79960
rect 145386 79908 145392 79960
rect 145788 79908 145794 79960
rect 145846 79908 145852 79960
rect 145880 79908 145886 79960
rect 145938 79908 145944 79960
rect 146064 79948 146070 79960
rect 146036 79908 146070 79948
rect 146122 79908 146128 79960
rect 146248 79948 146254 79960
rect 146220 79908 146254 79948
rect 146306 79948 146312 79960
rect 146306 79920 146353 79948
rect 146306 79908 146312 79920
rect 146524 79908 146530 79960
rect 146582 79908 146588 79960
rect 143506 79852 143902 79880
rect 143948 79840 143954 79892
rect 144006 79840 144012 79892
rect 143856 79812 143862 79824
rect 143828 79772 143862 79812
rect 143914 79772 143920 79824
rect 143046 79716 143304 79744
rect 143414 79716 143448 79756
rect 141878 79636 141884 79688
rect 141936 79636 141942 79688
rect 141970 79636 141976 79688
rect 142028 79636 142034 79688
rect 142246 79636 142252 79688
rect 142304 79636 142310 79688
rect 141292 79512 141694 79540
rect 141292 79500 141298 79512
rect 142154 79472 142160 79484
rect 128326 79444 142160 79472
rect 142154 79432 142160 79444
rect 142212 79432 142218 79484
rect 142632 79472 142660 79704
rect 142706 79568 142712 79620
rect 142764 79608 142770 79620
rect 143074 79608 143080 79620
rect 142764 79580 143080 79608
rect 142764 79568 142770 79580
rect 143074 79568 143080 79580
rect 143132 79568 143138 79620
rect 143276 79552 143304 79716
rect 143442 79704 143448 79716
rect 143500 79704 143506 79756
rect 143534 79704 143540 79756
rect 143592 79704 143598 79756
rect 143350 79636 143356 79688
rect 143408 79676 143414 79688
rect 143552 79676 143580 79704
rect 143408 79648 143580 79676
rect 143408 79636 143414 79648
rect 143828 79552 143856 79772
rect 143966 79688 143994 79840
rect 143902 79636 143908 79688
rect 143960 79648 143994 79688
rect 143960 79636 143966 79648
rect 144104 79620 144132 79908
rect 144242 79880 144270 79908
rect 144196 79852 144270 79880
rect 144196 79824 144224 79852
rect 144592 79840 144598 79892
rect 144650 79840 144656 79892
rect 144868 79840 144874 79892
rect 144926 79840 144932 79892
rect 144178 79772 144184 79824
rect 144236 79772 144242 79824
rect 144316 79812 144322 79824
rect 144288 79772 144322 79812
rect 144374 79772 144380 79824
rect 144408 79772 144414 79824
rect 144466 79772 144472 79824
rect 144500 79772 144506 79824
rect 144558 79772 144564 79824
rect 144288 79620 144316 79772
rect 144086 79568 144092 79620
rect 144144 79568 144150 79620
rect 144270 79568 144276 79620
rect 144328 79568 144334 79620
rect 143258 79500 143264 79552
rect 143316 79500 143322 79552
rect 143810 79500 143816 79552
rect 143868 79500 143874 79552
rect 143074 79472 143080 79484
rect 142632 79444 143080 79472
rect 143074 79432 143080 79444
rect 143132 79432 143138 79484
rect 143718 79432 143724 79484
rect 143776 79472 143782 79484
rect 144426 79472 144454 79772
rect 143776 79444 144454 79472
rect 144518 79484 144546 79772
rect 144610 79552 144638 79840
rect 144730 79636 144736 79688
rect 144788 79676 144794 79688
rect 144886 79676 144914 79840
rect 144788 79648 144914 79676
rect 144788 79636 144794 79648
rect 144822 79568 144828 79620
rect 144880 79608 144886 79620
rect 145346 79608 145374 79908
rect 145420 79840 145426 79892
rect 145478 79880 145484 79892
rect 145696 79880 145702 79892
rect 145478 79840 145512 79880
rect 145484 79688 145512 79840
rect 145668 79840 145702 79880
rect 145754 79840 145760 79892
rect 145668 79688 145696 79840
rect 145806 79812 145834 79908
rect 145760 79784 145834 79812
rect 145760 79756 145788 79784
rect 145898 79756 145926 79908
rect 145742 79704 145748 79756
rect 145800 79704 145806 79756
rect 145834 79704 145840 79756
rect 145892 79716 145926 79756
rect 145892 79704 145898 79716
rect 146036 79688 146064 79908
rect 145466 79636 145472 79688
rect 145524 79636 145530 79688
rect 145650 79636 145656 79688
rect 145708 79636 145714 79688
rect 146018 79636 146024 79688
rect 146076 79636 146082 79688
rect 146110 79636 146116 79688
rect 146168 79676 146174 79688
rect 146220 79676 146248 79908
rect 146340 79880 146346 79892
rect 146312 79840 146346 79880
rect 146398 79840 146404 79892
rect 146432 79840 146438 79892
rect 146490 79840 146496 79892
rect 146312 79756 146340 79840
rect 146450 79756 146478 79840
rect 146294 79704 146300 79756
rect 146352 79704 146358 79756
rect 146386 79704 146392 79756
rect 146444 79716 146478 79756
rect 146542 79756 146570 79908
rect 146542 79716 146576 79756
rect 146444 79704 146450 79716
rect 146570 79704 146576 79716
rect 146628 79704 146634 79756
rect 146680 79688 146708 79988
rect 147002 79960 147030 79988
rect 146800 79908 146806 79960
rect 146858 79948 146864 79960
rect 146858 79908 146892 79948
rect 146984 79908 146990 79960
rect 147042 79908 147048 79960
rect 147076 79908 147082 79960
rect 147134 79908 147140 79960
rect 147168 79908 147174 79960
rect 147226 79908 147232 79960
rect 147352 79908 147358 79960
rect 147410 79908 147416 79960
rect 147812 79948 147818 79960
rect 147784 79908 147818 79948
rect 147870 79908 147876 79960
rect 147996 79948 148002 79960
rect 147968 79908 148002 79948
rect 148054 79908 148060 79960
rect 148088 79908 148094 79960
rect 148146 79908 148152 79960
rect 148180 79908 148186 79960
rect 148238 79908 148244 79960
rect 148732 79908 148738 79960
rect 148790 79908 148796 79960
rect 146864 79688 146892 79908
rect 147094 79824 147122 79908
rect 147030 79772 147036 79824
rect 147088 79784 147122 79824
rect 147186 79824 147214 79908
rect 147370 79824 147398 79908
rect 147444 79840 147450 79892
rect 147502 79840 147508 79892
rect 147186 79784 147220 79824
rect 147088 79772 147094 79784
rect 147214 79772 147220 79784
rect 147272 79772 147278 79824
rect 147306 79772 147312 79824
rect 147364 79784 147398 79824
rect 147364 79772 147370 79784
rect 147462 79756 147490 79840
rect 147398 79704 147404 79756
rect 147456 79716 147490 79756
rect 147456 79704 147462 79716
rect 146168 79648 146248 79676
rect 146168 79636 146174 79648
rect 146662 79636 146668 79688
rect 146720 79636 146726 79688
rect 146846 79636 146852 79688
rect 146904 79636 146910 79688
rect 144880 79580 145374 79608
rect 144880 79568 144886 79580
rect 144610 79512 144644 79552
rect 144638 79500 144644 79512
rect 144696 79500 144702 79552
rect 144518 79444 144552 79484
rect 143776 79432 143782 79444
rect 144546 79432 144552 79444
rect 144604 79432 144610 79484
rect 147122 79432 147128 79484
rect 147180 79472 147186 79484
rect 147784 79472 147812 79908
rect 147968 79688 147996 79908
rect 148106 79756 148134 79908
rect 148042 79704 148048 79756
rect 148100 79716 148134 79756
rect 148100 79704 148106 79716
rect 148198 79688 148226 79908
rect 148272 79840 148278 79892
rect 148330 79840 148336 79892
rect 148364 79840 148370 79892
rect 148422 79880 148428 79892
rect 148422 79840 148456 79880
rect 148548 79840 148554 79892
rect 148606 79880 148612 79892
rect 148606 79840 148640 79880
rect 147950 79636 147956 79688
rect 148008 79636 148014 79688
rect 148134 79636 148140 79688
rect 148192 79648 148226 79688
rect 148290 79688 148318 79840
rect 148290 79648 148324 79688
rect 148192 79636 148198 79648
rect 148318 79636 148324 79648
rect 148376 79636 148382 79688
rect 148428 79676 148456 79840
rect 148612 79756 148640 79840
rect 148750 79824 148778 79908
rect 148842 79892 148870 80532
rect 149210 80016 149238 80600
rect 151786 80288 151814 80940
rect 158686 80900 158714 81008
rect 156064 80872 158714 80900
rect 156064 80356 156092 80872
rect 150682 80260 151814 80288
rect 152062 80328 156092 80356
rect 156984 80804 158714 80832
rect 149210 79988 150434 80016
rect 149210 79960 149238 79988
rect 149192 79908 149198 79960
rect 149250 79908 149256 79960
rect 149836 79908 149842 79960
rect 149894 79908 149900 79960
rect 150112 79908 150118 79960
rect 150170 79948 150176 79960
rect 150170 79908 150204 79948
rect 150296 79908 150302 79960
rect 150354 79908 150360 79960
rect 148824 79840 148830 79892
rect 148882 79840 148888 79892
rect 149284 79840 149290 79892
rect 149342 79840 149348 79892
rect 149376 79840 149382 79892
rect 149434 79880 149440 79892
rect 149434 79840 149468 79880
rect 148686 79772 148692 79824
rect 148744 79784 148778 79824
rect 148744 79772 148750 79784
rect 148594 79704 148600 79756
rect 148652 79704 148658 79756
rect 148842 79744 148870 79840
rect 149302 79812 149330 79840
rect 149302 79784 149376 79812
rect 149238 79744 149244 79756
rect 148842 79716 149244 79744
rect 149238 79704 149244 79716
rect 149296 79704 149302 79756
rect 148428 79648 148824 79676
rect 147858 79568 147864 79620
rect 147916 79608 147922 79620
rect 148686 79608 148692 79620
rect 147916 79580 148692 79608
rect 147916 79568 147922 79580
rect 148686 79568 148692 79580
rect 148744 79568 148750 79620
rect 148502 79500 148508 79552
rect 148560 79540 148566 79552
rect 148796 79540 148824 79648
rect 148560 79512 148824 79540
rect 148560 79500 148566 79512
rect 148870 79472 148876 79484
rect 147180 79444 148876 79472
rect 147180 79432 147186 79444
rect 148870 79432 148876 79444
rect 148928 79432 148934 79484
rect 111150 79364 111156 79416
rect 111208 79404 111214 79416
rect 131758 79404 131764 79416
rect 111208 79376 131764 79404
rect 111208 79364 111214 79376
rect 131758 79364 131764 79376
rect 131816 79364 131822 79416
rect 131850 79364 131856 79416
rect 131908 79404 131914 79416
rect 142982 79404 142988 79416
rect 131908 79376 142988 79404
rect 131908 79364 131914 79376
rect 142982 79364 142988 79376
rect 143040 79364 143046 79416
rect 149348 79404 149376 79784
rect 149440 79472 149468 79840
rect 149854 79540 149882 79908
rect 150020 79840 150026 79892
rect 150078 79880 150084 79892
rect 150078 79840 150112 79880
rect 150084 79608 150112 79840
rect 150176 79688 150204 79908
rect 150314 79824 150342 79908
rect 150250 79772 150256 79824
rect 150308 79784 150342 79824
rect 150308 79772 150314 79784
rect 150406 79756 150434 79988
rect 150682 79960 150710 80260
rect 150958 79988 151998 80016
rect 150958 79960 150986 79988
rect 150664 79908 150670 79960
rect 150722 79908 150728 79960
rect 150940 79908 150946 79960
rect 150998 79908 151004 79960
rect 151400 79948 151406 79960
rect 151234 79920 151406 79948
rect 151124 79840 151130 79892
rect 151182 79840 151188 79892
rect 151142 79812 151170 79840
rect 150342 79704 150348 79756
rect 150400 79716 150434 79756
rect 150728 79784 151170 79812
rect 150400 79704 150406 79716
rect 150158 79636 150164 79688
rect 150216 79636 150222 79688
rect 150728 79620 150756 79784
rect 151234 79744 151262 79920
rect 151400 79908 151406 79920
rect 151458 79908 151464 79960
rect 151492 79880 151498 79892
rect 151464 79840 151498 79880
rect 151550 79840 151556 79892
rect 151970 79880 151998 79988
rect 152062 79960 152090 80328
rect 156984 80288 157012 80804
rect 158686 80628 158714 80804
rect 159146 80764 159174 81008
rect 182008 81008 186780 81036
rect 182008 80968 182036 81008
rect 186774 80996 186780 81008
rect 186832 80996 186838 81048
rect 200758 80968 200764 80980
rect 171152 80940 182036 80968
rect 182146 80940 200764 80968
rect 171152 80764 171180 80940
rect 182146 80900 182174 80940
rect 200758 80928 200764 80940
rect 200816 80928 200822 80980
rect 159146 80736 171180 80764
rect 178604 80872 182174 80900
rect 159054 80668 170996 80696
rect 159054 80628 159082 80668
rect 158686 80600 159082 80628
rect 170968 80628 170996 80668
rect 178604 80628 178632 80872
rect 187418 80860 187424 80912
rect 187476 80900 187482 80912
rect 206186 80900 206192 80912
rect 187476 80872 206192 80900
rect 187476 80860 187482 80872
rect 206186 80860 206192 80872
rect 206244 80900 206250 80912
rect 234614 80900 234620 80912
rect 206244 80872 234620 80900
rect 206244 80860 206250 80872
rect 234614 80860 234620 80872
rect 234672 80860 234678 80912
rect 186774 80792 186780 80844
rect 186832 80832 186838 80844
rect 252554 80832 252560 80844
rect 186832 80804 252560 80832
rect 186832 80792 186838 80804
rect 252554 80792 252560 80804
rect 252612 80792 252618 80844
rect 188154 80764 188160 80776
rect 178880 80736 188160 80764
rect 178770 80628 178776 80640
rect 170968 80600 171088 80628
rect 178604 80600 178776 80628
rect 171060 80560 171088 80600
rect 178770 80588 178776 80600
rect 178828 80588 178834 80640
rect 178880 80560 178908 80736
rect 188154 80724 188160 80736
rect 188212 80764 188218 80776
rect 270494 80764 270500 80776
rect 188212 80736 270500 80764
rect 188212 80724 188218 80736
rect 270494 80724 270500 80736
rect 270552 80724 270558 80776
rect 195146 80696 195152 80708
rect 182146 80668 195152 80696
rect 182146 80628 182174 80668
rect 195146 80656 195152 80668
rect 195204 80696 195210 80708
rect 358814 80696 358820 80708
rect 195204 80668 358820 80696
rect 195204 80656 195210 80668
rect 358814 80656 358820 80668
rect 358872 80656 358878 80708
rect 171060 80532 178908 80560
rect 179386 80600 182174 80628
rect 177758 80452 177764 80504
rect 177816 80492 177822 80504
rect 179386 80492 179414 80600
rect 177816 80464 179414 80492
rect 177816 80452 177822 80464
rect 179598 80424 179604 80436
rect 173222 80396 179604 80424
rect 173222 80356 173250 80396
rect 179598 80384 179604 80396
rect 179656 80424 179662 80436
rect 179656 80396 183554 80424
rect 179656 80384 179662 80396
rect 178034 80356 178040 80368
rect 154316 80260 157012 80288
rect 158686 80328 173250 80356
rect 173314 80328 178040 80356
rect 152614 79988 153378 80016
rect 152044 79908 152050 79960
rect 152102 79908 152108 79960
rect 152614 79880 152642 79988
rect 153056 79948 153062 79960
rect 153028 79908 153062 79948
rect 153114 79908 153120 79960
rect 153148 79908 153154 79960
rect 153206 79908 153212 79960
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 151970 79852 152642 79880
rect 152688 79840 152694 79892
rect 152746 79880 152752 79892
rect 152746 79852 152964 79880
rect 152746 79840 152752 79852
rect 151308 79772 151314 79824
rect 151366 79772 151372 79824
rect 150912 79716 151262 79744
rect 150526 79608 150532 79620
rect 150084 79580 150532 79608
rect 150526 79568 150532 79580
rect 150584 79568 150590 79620
rect 150710 79568 150716 79620
rect 150768 79568 150774 79620
rect 150912 79608 150940 79716
rect 151326 79688 151354 79772
rect 151464 79756 151492 79840
rect 151446 79704 151452 79756
rect 151504 79704 151510 79756
rect 151326 79648 151360 79688
rect 151354 79636 151360 79648
rect 151412 79636 151418 79688
rect 151262 79608 151268 79620
rect 150912 79580 151268 79608
rect 150912 79552 150940 79580
rect 151262 79568 151268 79580
rect 151320 79568 151326 79620
rect 152550 79608 152556 79620
rect 152292 79580 152556 79608
rect 152292 79552 152320 79580
rect 152550 79568 152556 79580
rect 152608 79568 152614 79620
rect 149854 79512 150112 79540
rect 149974 79472 149980 79484
rect 149440 79444 149980 79472
rect 149974 79432 149980 79444
rect 150032 79432 150038 79484
rect 149698 79404 149704 79416
rect 149348 79376 149704 79404
rect 149698 79364 149704 79376
rect 149756 79364 149762 79416
rect 149882 79364 149888 79416
rect 149940 79404 149946 79416
rect 150084 79404 150112 79512
rect 150894 79500 150900 79552
rect 150952 79500 150958 79552
rect 152274 79500 152280 79552
rect 152332 79500 152338 79552
rect 150802 79432 150808 79484
rect 150860 79472 150866 79484
rect 151538 79472 151544 79484
rect 150860 79444 151544 79472
rect 150860 79432 150866 79444
rect 151538 79432 151544 79444
rect 151596 79432 151602 79484
rect 151722 79432 151728 79484
rect 151780 79472 151786 79484
rect 151780 79444 151952 79472
rect 151780 79432 151786 79444
rect 149940 79376 150112 79404
rect 149940 79364 149946 79376
rect 104894 79296 104900 79348
rect 104952 79336 104958 79348
rect 105998 79336 106004 79348
rect 104952 79308 106004 79336
rect 104952 79296 104958 79308
rect 105998 79296 106004 79308
rect 106056 79296 106062 79348
rect 109770 79296 109776 79348
rect 109828 79336 109834 79348
rect 132310 79336 132316 79348
rect 109828 79308 132316 79336
rect 109828 79296 109834 79308
rect 132310 79296 132316 79308
rect 132368 79296 132374 79348
rect 133230 79296 133236 79348
rect 133288 79336 133294 79348
rect 135530 79336 135536 79348
rect 133288 79308 135536 79336
rect 133288 79296 133294 79308
rect 135530 79296 135536 79308
rect 135588 79296 135594 79348
rect 138290 79296 138296 79348
rect 138348 79336 138354 79348
rect 138934 79336 138940 79348
rect 138348 79308 138940 79336
rect 138348 79296 138354 79308
rect 138934 79296 138940 79308
rect 138992 79296 138998 79348
rect 149238 79336 149244 79348
rect 142126 79308 149244 79336
rect 123662 79228 123668 79280
rect 123720 79268 123726 79280
rect 142126 79268 142154 79308
rect 149238 79296 149244 79308
rect 149296 79296 149302 79348
rect 147950 79268 147956 79280
rect 123720 79240 142154 79268
rect 142908 79240 147956 79268
rect 123720 79228 123726 79240
rect 119338 79160 119344 79212
rect 119396 79200 119402 79212
rect 141326 79200 141332 79212
rect 119396 79172 141332 79200
rect 119396 79160 119402 79172
rect 141326 79160 141332 79172
rect 141384 79160 141390 79212
rect 142908 79200 142936 79240
rect 147950 79228 147956 79240
rect 148008 79228 148014 79280
rect 151446 79228 151452 79280
rect 151504 79268 151510 79280
rect 151924 79268 151952 79444
rect 152090 79432 152096 79484
rect 152148 79472 152154 79484
rect 152826 79472 152832 79484
rect 152148 79444 152832 79472
rect 152148 79432 152154 79444
rect 152826 79432 152832 79444
rect 152884 79432 152890 79484
rect 152642 79364 152648 79416
rect 152700 79404 152706 79416
rect 152936 79404 152964 79852
rect 152700 79376 152964 79404
rect 152700 79364 152706 79376
rect 152182 79296 152188 79348
rect 152240 79336 152246 79348
rect 153028 79336 153056 79908
rect 153166 79824 153194 79908
rect 153102 79772 153108 79824
rect 153160 79784 153194 79824
rect 153160 79772 153166 79784
rect 153258 79756 153286 79908
rect 153194 79704 153200 79756
rect 153252 79716 153286 79756
rect 153252 79704 153258 79716
rect 153350 79608 153378 79988
rect 153424 79908 153430 79960
rect 153482 79948 153488 79960
rect 154316 79948 154344 80260
rect 158686 80220 158714 80328
rect 173314 80288 173342 80328
rect 178034 80316 178040 80328
rect 178092 80316 178098 80368
rect 179874 80288 179880 80300
rect 153482 79920 154344 79948
rect 154408 80192 158714 80220
rect 173222 80260 173342 80288
rect 174188 80260 179880 80288
rect 153482 79908 153488 79920
rect 153700 79840 153706 79892
rect 153758 79840 153764 79892
rect 154068 79840 154074 79892
rect 154126 79840 154132 79892
rect 154160 79840 154166 79892
rect 154218 79880 154224 79892
rect 154218 79852 154344 79880
rect 154218 79840 154224 79852
rect 153718 79744 153746 79840
rect 154086 79756 154114 79840
rect 153718 79716 153976 79744
rect 154086 79716 154120 79756
rect 153948 79688 153976 79716
rect 154114 79704 154120 79716
rect 154172 79704 154178 79756
rect 154316 79688 154344 79852
rect 153930 79636 153936 79688
rect 153988 79636 153994 79688
rect 154298 79636 154304 79688
rect 154356 79636 154362 79688
rect 154408 79608 154436 80192
rect 166506 80056 171502 80084
rect 163746 79988 165706 80016
rect 163746 79960 163774 79988
rect 154528 79908 154534 79960
rect 154586 79908 154592 79960
rect 154620 79908 154626 79960
rect 154678 79908 154684 79960
rect 154712 79908 154718 79960
rect 154770 79948 154776 79960
rect 155172 79948 155178 79960
rect 154770 79920 155080 79948
rect 154770 79908 154776 79920
rect 154546 79688 154574 79908
rect 154638 79756 154666 79908
rect 154638 79716 154672 79756
rect 154666 79704 154672 79716
rect 154724 79704 154730 79756
rect 155052 79688 155080 79920
rect 155144 79908 155178 79948
rect 155230 79908 155236 79960
rect 155264 79908 155270 79960
rect 155322 79908 155328 79960
rect 155724 79908 155730 79960
rect 155782 79908 155788 79960
rect 155908 79908 155914 79960
rect 155966 79908 155972 79960
rect 156092 79908 156098 79960
rect 156150 79908 156156 79960
rect 156276 79908 156282 79960
rect 156334 79908 156340 79960
rect 156460 79908 156466 79960
rect 156518 79908 156524 79960
rect 156552 79908 156558 79960
rect 156610 79908 156616 79960
rect 156828 79908 156834 79960
rect 156886 79908 156892 79960
rect 156920 79908 156926 79960
rect 156978 79908 156984 79960
rect 157288 79908 157294 79960
rect 157346 79908 157352 79960
rect 157656 79908 157662 79960
rect 157714 79908 157720 79960
rect 158300 79948 158306 79960
rect 157812 79920 158306 79948
rect 154482 79636 154488 79688
rect 154540 79648 154574 79688
rect 154540 79636 154546 79648
rect 155034 79636 155040 79688
rect 155092 79636 155098 79688
rect 153350 79580 154436 79608
rect 152240 79308 153056 79336
rect 153166 79512 154574 79540
rect 152240 79296 152246 79308
rect 151504 79240 151952 79268
rect 151504 79228 151510 79240
rect 141896 79172 142936 79200
rect 120626 79092 120632 79144
rect 120684 79132 120690 79144
rect 141896 79132 141924 79172
rect 142982 79160 142988 79212
rect 143040 79200 143046 79212
rect 153166 79200 153194 79512
rect 154546 79268 154574 79512
rect 155144 79472 155172 79908
rect 155282 79824 155310 79908
rect 155264 79772 155270 79824
rect 155322 79772 155328 79824
rect 155632 79772 155638 79824
rect 155690 79772 155696 79824
rect 155218 79636 155224 79688
rect 155276 79676 155282 79688
rect 155650 79676 155678 79772
rect 155276 79648 155678 79676
rect 155276 79636 155282 79648
rect 155742 79620 155770 79908
rect 155678 79568 155684 79620
rect 155736 79580 155770 79620
rect 155736 79568 155742 79580
rect 155310 79472 155316 79484
rect 155144 79444 155316 79472
rect 155310 79432 155316 79444
rect 155368 79432 155374 79484
rect 155926 79472 155954 79908
rect 156110 79540 156138 79908
rect 156294 79824 156322 79908
rect 156276 79772 156282 79824
rect 156334 79772 156340 79824
rect 156478 79744 156506 79908
rect 156570 79812 156598 79908
rect 156570 79784 156736 79812
rect 156478 79716 156552 79744
rect 156524 79620 156552 79716
rect 156708 79620 156736 79784
rect 156506 79568 156512 79620
rect 156564 79568 156570 79620
rect 156690 79568 156696 79620
rect 156748 79568 156754 79620
rect 156322 79540 156328 79552
rect 156110 79512 156328 79540
rect 156322 79500 156328 79512
rect 156380 79500 156386 79552
rect 156414 79472 156420 79484
rect 155926 79444 156420 79472
rect 156414 79432 156420 79444
rect 156472 79432 156478 79484
rect 156046 79364 156052 79416
rect 156104 79404 156110 79416
rect 156846 79404 156874 79908
rect 156938 79824 156966 79908
rect 156938 79784 156972 79824
rect 156966 79772 156972 79784
rect 157024 79772 157030 79824
rect 156966 79500 156972 79552
rect 157024 79540 157030 79552
rect 157306 79540 157334 79908
rect 157674 79880 157702 79908
rect 157024 79512 157334 79540
rect 157490 79852 157702 79880
rect 157024 79500 157030 79512
rect 157490 79484 157518 79852
rect 157564 79772 157570 79824
rect 157622 79772 157628 79824
rect 157582 79552 157610 79772
rect 157582 79512 157616 79552
rect 157610 79500 157616 79512
rect 157668 79500 157674 79552
rect 157812 79484 157840 79920
rect 158300 79908 158306 79920
rect 158358 79908 158364 79960
rect 159036 79908 159042 79960
rect 159094 79908 159100 79960
rect 159128 79908 159134 79960
rect 159186 79908 159192 79960
rect 159588 79908 159594 79960
rect 159646 79908 159652 79960
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160508 79908 160514 79960
rect 160566 79908 160572 79960
rect 160876 79908 160882 79960
rect 160934 79908 160940 79960
rect 161060 79908 161066 79960
rect 161118 79908 161124 79960
rect 161152 79908 161158 79960
rect 161210 79908 161216 79960
rect 161244 79908 161250 79960
rect 161302 79948 161308 79960
rect 161302 79920 161474 79948
rect 161302 79908 161308 79920
rect 158208 79840 158214 79892
rect 158266 79880 158272 79892
rect 158266 79852 158392 79880
rect 158266 79840 158272 79852
rect 158024 79772 158030 79824
rect 158082 79772 158088 79824
rect 158042 79688 158070 79772
rect 158364 79688 158392 79852
rect 158484 79840 158490 79892
rect 158542 79880 158548 79892
rect 158668 79880 158674 79892
rect 158542 79840 158576 79880
rect 158042 79648 158076 79688
rect 158070 79636 158076 79648
rect 158128 79636 158134 79688
rect 158346 79636 158352 79688
rect 158404 79636 158410 79688
rect 158548 79620 158576 79840
rect 158640 79840 158674 79880
rect 158726 79840 158732 79892
rect 158760 79840 158766 79892
rect 158818 79840 158824 79892
rect 158640 79620 158668 79840
rect 158530 79568 158536 79620
rect 158588 79568 158594 79620
rect 158622 79568 158628 79620
rect 158680 79568 158686 79620
rect 157490 79444 157524 79484
rect 157518 79432 157524 79444
rect 157576 79432 157582 79484
rect 157794 79432 157800 79484
rect 157852 79432 157858 79484
rect 156104 79376 156874 79404
rect 158778 79404 158806 79840
rect 158898 79500 158904 79552
rect 158956 79540 158962 79552
rect 159054 79540 159082 79908
rect 158956 79512 159082 79540
rect 158956 79500 158962 79512
rect 159146 79484 159174 79908
rect 159606 79824 159634 79908
rect 159772 79840 159778 79892
rect 159830 79840 159836 79892
rect 159542 79772 159548 79824
rect 159600 79784 159634 79824
rect 159600 79772 159606 79784
rect 159790 79744 159818 79840
rect 160434 79824 160462 79908
rect 160370 79772 160376 79824
rect 160428 79784 160462 79824
rect 160428 79772 160434 79784
rect 160526 79756 160554 79908
rect 160692 79880 160698 79892
rect 159376 79716 159818 79744
rect 159376 79484 159404 79716
rect 160462 79704 160468 79756
rect 160520 79716 160554 79756
rect 160664 79840 160698 79880
rect 160750 79840 160756 79892
rect 160784 79840 160790 79892
rect 160842 79840 160848 79892
rect 160520 79704 160526 79716
rect 160664 79620 160692 79840
rect 160802 79756 160830 79840
rect 160738 79704 160744 79756
rect 160796 79716 160830 79756
rect 160796 79704 160802 79716
rect 160894 79688 160922 79908
rect 161078 79812 161106 79908
rect 160830 79636 160836 79688
rect 160888 79648 160922 79688
rect 161032 79784 161106 79812
rect 160888 79636 160894 79648
rect 160646 79568 160652 79620
rect 160704 79568 160710 79620
rect 160922 79568 160928 79620
rect 160980 79608 160986 79620
rect 161032 79608 161060 79784
rect 161170 79756 161198 79908
rect 161336 79772 161342 79824
rect 161394 79772 161400 79824
rect 161106 79704 161112 79756
rect 161164 79716 161198 79756
rect 161164 79704 161170 79716
rect 161198 79636 161204 79688
rect 161256 79676 161262 79688
rect 161354 79676 161382 79772
rect 161256 79648 161382 79676
rect 161256 79636 161262 79648
rect 160980 79580 161060 79608
rect 160980 79568 160986 79580
rect 161290 79568 161296 79620
rect 161348 79608 161354 79620
rect 161446 79608 161474 79920
rect 161612 79908 161618 79960
rect 161670 79908 161676 79960
rect 161980 79908 161986 79960
rect 162038 79908 162044 79960
rect 162164 79908 162170 79960
rect 162222 79948 162228 79960
rect 162222 79908 162256 79948
rect 162992 79908 162998 79960
rect 163050 79908 163056 79960
rect 163084 79908 163090 79960
rect 163142 79908 163148 79960
rect 163360 79908 163366 79960
rect 163418 79908 163424 79960
rect 163728 79908 163734 79960
rect 163786 79908 163792 79960
rect 164004 79908 164010 79960
rect 164062 79908 164068 79960
rect 164096 79908 164102 79960
rect 164154 79908 164160 79960
rect 164464 79908 164470 79960
rect 164522 79908 164528 79960
rect 164832 79908 164838 79960
rect 164890 79908 164896 79960
rect 164924 79908 164930 79960
rect 164982 79908 164988 79960
rect 165200 79908 165206 79960
rect 165258 79908 165264 79960
rect 161630 79824 161658 79908
rect 161630 79784 161664 79824
rect 161658 79772 161664 79784
rect 161716 79772 161722 79824
rect 161888 79812 161894 79824
rect 161768 79784 161894 79812
rect 161348 79580 161474 79608
rect 161768 79608 161796 79784
rect 161888 79772 161894 79784
rect 161946 79772 161952 79824
rect 161998 79744 162026 79908
rect 161860 79716 162026 79744
rect 161860 79688 161888 79716
rect 162228 79688 162256 79908
rect 162348 79840 162354 79892
rect 162406 79840 162412 79892
rect 162532 79840 162538 79892
rect 162590 79840 162596 79892
rect 162624 79840 162630 79892
rect 162682 79880 162688 79892
rect 162682 79840 162716 79880
rect 162808 79840 162814 79892
rect 162866 79840 162872 79892
rect 163010 79880 163038 79908
rect 162964 79852 163038 79880
rect 161842 79636 161848 79688
rect 161900 79636 161906 79688
rect 162210 79636 162216 79688
rect 162268 79636 162274 79688
rect 162366 79620 162394 79840
rect 162550 79756 162578 79840
rect 162688 79756 162716 79840
rect 162550 79716 162584 79756
rect 162578 79704 162584 79716
rect 162636 79704 162642 79756
rect 162670 79704 162676 79756
rect 162728 79704 162734 79756
rect 161934 79608 161940 79620
rect 161768 79580 161940 79608
rect 161348 79568 161354 79580
rect 161934 79568 161940 79580
rect 161992 79568 161998 79620
rect 162366 79580 162400 79620
rect 162394 79568 162400 79580
rect 162452 79568 162458 79620
rect 159634 79500 159640 79552
rect 159692 79540 159698 79552
rect 159910 79540 159916 79552
rect 159692 79512 159916 79540
rect 159692 79500 159698 79512
rect 159910 79500 159916 79512
rect 159968 79500 159974 79552
rect 159082 79432 159088 79484
rect 159140 79444 159174 79484
rect 159140 79432 159146 79444
rect 159358 79432 159364 79484
rect 159416 79432 159422 79484
rect 159726 79404 159732 79416
rect 158778 79376 159732 79404
rect 156104 79364 156110 79376
rect 159726 79364 159732 79376
rect 159784 79364 159790 79416
rect 161566 79364 161572 79416
rect 161624 79404 161630 79416
rect 162826 79404 162854 79840
rect 162964 79756 162992 79852
rect 163102 79812 163130 79908
rect 163268 79840 163274 79892
rect 163326 79840 163332 79892
rect 163056 79784 163130 79812
rect 162946 79704 162952 79756
rect 163004 79704 163010 79756
rect 163056 79620 163084 79784
rect 163176 79772 163182 79824
rect 163234 79772 163240 79824
rect 163194 79744 163222 79772
rect 163148 79716 163222 79744
rect 163038 79568 163044 79620
rect 163096 79568 163102 79620
rect 163148 79552 163176 79716
rect 163286 79688 163314 79840
rect 163222 79636 163228 79688
rect 163280 79648 163314 79688
rect 163280 79636 163286 79648
rect 163378 79620 163406 79908
rect 163820 79880 163826 79892
rect 163792 79840 163826 79880
rect 163878 79840 163884 79892
rect 163452 79772 163458 79824
rect 163510 79772 163516 79824
rect 163314 79568 163320 79620
rect 163372 79580 163406 79620
rect 163372 79568 163378 79580
rect 163130 79500 163136 79552
rect 163188 79500 163194 79552
rect 163470 79472 163498 79772
rect 163792 79620 163820 79840
rect 163774 79568 163780 79620
rect 163832 79568 163838 79620
rect 163866 79568 163872 79620
rect 163924 79608 163930 79620
rect 164022 79608 164050 79908
rect 164114 79824 164142 79908
rect 164188 79840 164194 79892
rect 164246 79840 164252 79892
rect 164280 79840 164286 79892
rect 164338 79880 164344 79892
rect 164338 79840 164372 79880
rect 164096 79772 164102 79824
rect 164154 79772 164160 79824
rect 163924 79580 164050 79608
rect 164206 79620 164234 79840
rect 164344 79756 164372 79840
rect 164326 79704 164332 79756
rect 164384 79704 164390 79756
rect 164206 79580 164240 79620
rect 163924 79568 163930 79580
rect 164234 79568 164240 79580
rect 164292 79568 164298 79620
rect 164482 79608 164510 79908
rect 164850 79744 164878 79908
rect 164942 79756 164970 79908
rect 165218 79824 165246 79908
rect 165476 79840 165482 79892
rect 165534 79840 165540 79892
rect 165218 79784 165252 79824
rect 165246 79772 165252 79784
rect 165304 79772 165310 79824
rect 164344 79580 164510 79608
rect 164712 79716 164878 79744
rect 164712 79608 164740 79716
rect 164924 79704 164930 79756
rect 164982 79704 164988 79756
rect 164786 79636 164792 79688
rect 164844 79676 164850 79688
rect 165494 79676 165522 79840
rect 164844 79648 165522 79676
rect 164844 79636 164850 79648
rect 165356 79620 165384 79648
rect 164878 79608 164884 79620
rect 164712 79580 164884 79608
rect 163590 79472 163596 79484
rect 163470 79444 163596 79472
rect 163590 79432 163596 79444
rect 163648 79432 163654 79484
rect 164344 79472 164372 79580
rect 164878 79568 164884 79580
rect 164936 79568 164942 79620
rect 165062 79608 165068 79620
rect 164988 79580 165068 79608
rect 164988 79552 165016 79580
rect 165062 79568 165068 79580
rect 165120 79568 165126 79620
rect 165338 79568 165344 79620
rect 165396 79568 165402 79620
rect 164418 79500 164424 79552
rect 164476 79540 164482 79552
rect 164694 79540 164700 79552
rect 164476 79512 164700 79540
rect 164476 79500 164482 79512
rect 164694 79500 164700 79512
rect 164752 79500 164758 79552
rect 164970 79500 164976 79552
rect 165028 79500 165034 79552
rect 165678 79540 165706 79988
rect 166506 79960 166534 80056
rect 165936 79908 165942 79960
rect 165994 79908 166000 79960
rect 166120 79908 166126 79960
rect 166178 79908 166184 79960
rect 166212 79908 166218 79960
rect 166270 79908 166276 79960
rect 166304 79908 166310 79960
rect 166362 79908 166368 79960
rect 166396 79908 166402 79960
rect 166454 79908 166460 79960
rect 166488 79908 166494 79960
rect 166546 79908 166552 79960
rect 165752 79772 165758 79824
rect 165810 79772 165816 79824
rect 165770 79688 165798 79772
rect 165770 79648 165804 79688
rect 165798 79636 165804 79648
rect 165856 79636 165862 79688
rect 165954 79608 165982 79908
rect 166138 79824 166166 79908
rect 166074 79772 166080 79824
rect 166132 79784 166166 79824
rect 166132 79772 166138 79784
rect 166230 79756 166258 79908
rect 166166 79704 166172 79756
rect 166224 79716 166258 79756
rect 166224 79704 166230 79716
rect 166322 79676 166350 79908
rect 166414 79756 166442 79908
rect 166764 79840 166770 79892
rect 166822 79840 166828 79892
rect 166856 79840 166862 79892
rect 166914 79840 166920 79892
rect 166414 79716 166448 79756
rect 166442 79704 166448 79716
rect 166500 79704 166506 79756
rect 166626 79676 166632 79688
rect 166322 79648 166632 79676
rect 166626 79636 166632 79648
rect 166684 79636 166690 79688
rect 166350 79608 166356 79620
rect 165954 79580 166356 79608
rect 166350 79568 166356 79580
rect 166408 79568 166414 79620
rect 166782 79552 166810 79840
rect 166874 79608 166902 79840
rect 166994 79608 167000 79620
rect 166874 79580 167000 79608
rect 166994 79568 167000 79580
rect 167052 79568 167058 79620
rect 165982 79540 165988 79552
rect 165678 79512 165988 79540
rect 165982 79500 165988 79512
rect 166040 79500 166046 79552
rect 166718 79500 166724 79552
rect 166776 79512 166810 79552
rect 166776 79500 166782 79512
rect 165062 79472 165068 79484
rect 164344 79444 165068 79472
rect 165062 79432 165068 79444
rect 165120 79432 165126 79484
rect 165614 79432 165620 79484
rect 165672 79472 165678 79484
rect 167104 79472 167132 80056
rect 170140 79988 170582 80016
rect 167224 79908 167230 79960
rect 167282 79908 167288 79960
rect 167684 79908 167690 79960
rect 167742 79948 167748 79960
rect 167742 79920 168052 79948
rect 167742 79908 167748 79920
rect 167242 79744 167270 79908
rect 167242 79716 167500 79744
rect 167178 79568 167184 79620
rect 167236 79608 167242 79620
rect 167472 79608 167500 79716
rect 167236 79580 167500 79608
rect 167236 79568 167242 79580
rect 168024 79552 168052 79920
rect 168328 79908 168334 79960
rect 168386 79908 168392 79960
rect 168420 79908 168426 79960
rect 168478 79908 168484 79960
rect 168512 79908 168518 79960
rect 168570 79908 168576 79960
rect 168880 79908 168886 79960
rect 168938 79908 168944 79960
rect 169064 79908 169070 79960
rect 169122 79948 169128 79960
rect 169122 79920 169294 79948
rect 169122 79908 169128 79920
rect 168346 79824 168374 79908
rect 168438 79824 168466 79908
rect 168282 79772 168288 79824
rect 168340 79784 168374 79824
rect 168340 79772 168346 79784
rect 168420 79772 168426 79824
rect 168478 79772 168484 79824
rect 168530 79620 168558 79908
rect 168604 79772 168610 79824
rect 168662 79772 168668 79824
rect 168622 79744 168650 79772
rect 168622 79716 168696 79744
rect 168668 79620 168696 79716
rect 168530 79580 168564 79620
rect 168558 79568 168564 79580
rect 168616 79568 168622 79620
rect 168650 79568 168656 79620
rect 168708 79568 168714 79620
rect 168898 79552 168926 79908
rect 168972 79840 168978 79892
rect 169030 79840 169036 79892
rect 168990 79812 169018 79840
rect 169110 79812 169116 79824
rect 168990 79784 169116 79812
rect 169110 79772 169116 79784
rect 169168 79772 169174 79824
rect 169266 79620 169294 79920
rect 169708 79908 169714 79960
rect 169766 79908 169772 79960
rect 169800 79908 169806 79960
rect 169858 79908 169864 79960
rect 169984 79908 169990 79960
rect 170042 79948 170048 79960
rect 170042 79908 170076 79948
rect 169340 79840 169346 79892
rect 169398 79840 169404 79892
rect 169616 79880 169622 79892
rect 169588 79840 169622 79880
rect 169674 79840 169680 79892
rect 169202 79568 169208 79620
rect 169260 79580 169294 79620
rect 169358 79620 169386 79840
rect 169358 79580 169392 79620
rect 169260 79568 169266 79580
rect 169386 79568 169392 79580
rect 169444 79568 169450 79620
rect 168006 79500 168012 79552
rect 168064 79500 168070 79552
rect 168834 79500 168840 79552
rect 168892 79512 168926 79552
rect 169588 79540 169616 79840
rect 169726 79620 169754 79908
rect 169818 79756 169846 79908
rect 169892 79840 169898 79892
rect 169950 79880 169956 79892
rect 169950 79840 169984 79880
rect 169818 79716 169852 79756
rect 169846 79704 169852 79716
rect 169904 79704 169910 79756
rect 169662 79568 169668 79620
rect 169720 79580 169754 79620
rect 169720 79568 169726 79580
rect 169754 79540 169760 79552
rect 169588 79512 169760 79540
rect 168892 79500 168898 79512
rect 169754 79500 169760 79512
rect 169812 79500 169818 79552
rect 165672 79444 167132 79472
rect 165672 79432 165678 79444
rect 169386 79432 169392 79484
rect 169444 79472 169450 79484
rect 169956 79472 169984 79840
rect 170048 79688 170076 79908
rect 170030 79636 170036 79688
rect 170088 79636 170094 79688
rect 170140 79540 170168 79988
rect 170554 79960 170582 79988
rect 170260 79908 170266 79960
rect 170318 79948 170324 79960
rect 170318 79920 170490 79948
rect 170318 79908 170324 79920
rect 170352 79840 170358 79892
rect 170410 79840 170416 79892
rect 170370 79744 170398 79840
rect 170462 79812 170490 79920
rect 170536 79908 170542 79960
rect 170594 79908 170600 79960
rect 170720 79908 170726 79960
rect 170778 79908 170784 79960
rect 171088 79948 171094 79960
rect 171060 79908 171094 79948
rect 171146 79908 171152 79960
rect 171180 79908 171186 79960
rect 171238 79948 171244 79960
rect 171364 79948 171370 79960
rect 171238 79908 171272 79948
rect 170738 79812 170766 79908
rect 170904 79840 170910 79892
rect 170962 79880 170968 79892
rect 170962 79840 170996 79880
rect 170462 79784 170628 79812
rect 170738 79784 170904 79812
rect 170370 79716 170536 79744
rect 170214 79568 170220 79620
rect 170272 79608 170278 79620
rect 170508 79608 170536 79716
rect 170272 79580 170536 79608
rect 170272 79568 170278 79580
rect 170306 79540 170312 79552
rect 170140 79512 170312 79540
rect 170306 79500 170312 79512
rect 170364 79500 170370 79552
rect 170398 79500 170404 79552
rect 170456 79540 170462 79552
rect 170600 79540 170628 79784
rect 170876 79688 170904 79784
rect 170858 79636 170864 79688
rect 170916 79636 170922 79688
rect 170968 79608 170996 79840
rect 171060 79688 171088 79908
rect 171244 79756 171272 79908
rect 171336 79908 171370 79948
rect 171422 79908 171428 79960
rect 171336 79824 171364 79908
rect 171318 79772 171324 79824
rect 171376 79772 171382 79824
rect 171226 79704 171232 79756
rect 171284 79704 171290 79756
rect 171474 79744 171502 80056
rect 173222 80016 173250 80260
rect 174188 80152 174216 80260
rect 179874 80248 179880 80260
rect 179932 80248 179938 80300
rect 179322 80220 179328 80232
rect 171750 79988 173250 80016
rect 173314 80124 174216 80152
rect 174280 80192 179328 80220
rect 171750 79960 171778 79988
rect 173314 79960 173342 80124
rect 174280 80084 174308 80192
rect 179322 80180 179328 80192
rect 179380 80180 179386 80232
rect 178494 80152 178500 80164
rect 173498 80056 174308 80084
rect 174418 80124 178500 80152
rect 171732 79908 171738 79960
rect 171790 79908 171796 79960
rect 172008 79908 172014 79960
rect 172066 79908 172072 79960
rect 172376 79908 172382 79960
rect 172434 79908 172440 79960
rect 172836 79908 172842 79960
rect 172894 79908 172900 79960
rect 172928 79908 172934 79960
rect 172986 79908 172992 79960
rect 173020 79908 173026 79960
rect 173078 79948 173084 79960
rect 173078 79908 173112 79948
rect 173204 79908 173210 79960
rect 173262 79908 173268 79960
rect 173296 79908 173302 79960
rect 173354 79908 173360 79960
rect 173388 79908 173394 79960
rect 173446 79908 173452 79960
rect 171336 79716 171502 79744
rect 171042 79636 171048 79688
rect 171100 79636 171106 79688
rect 171134 79608 171140 79620
rect 170968 79580 171140 79608
rect 171134 79568 171140 79580
rect 171192 79568 171198 79620
rect 171336 79608 171364 79716
rect 171410 79636 171416 79688
rect 171468 79676 171474 79688
rect 171750 79676 171778 79908
rect 172026 79824 172054 79908
rect 172394 79824 172422 79908
rect 172026 79784 172060 79824
rect 172054 79772 172060 79784
rect 172112 79772 172118 79824
rect 172330 79772 172336 79824
rect 172388 79784 172422 79824
rect 172388 79772 172394 79784
rect 172854 79756 172882 79908
rect 172946 79824 172974 79908
rect 172946 79784 172980 79824
rect 172974 79772 172980 79784
rect 173032 79772 173038 79824
rect 172790 79704 172796 79756
rect 172848 79716 172882 79756
rect 173084 79744 173112 79908
rect 173222 79824 173250 79908
rect 173406 79824 173434 79908
rect 173222 79784 173256 79824
rect 173250 79772 173256 79784
rect 173308 79772 173314 79824
rect 173342 79772 173348 79824
rect 173400 79784 173434 79824
rect 173400 79772 173406 79784
rect 173498 79744 173526 80056
rect 173682 79988 173894 80016
rect 173682 79960 173710 79988
rect 173664 79908 173670 79960
rect 173722 79908 173728 79960
rect 173756 79908 173762 79960
rect 173814 79908 173820 79960
rect 173572 79840 173578 79892
rect 173630 79840 173636 79892
rect 173084 79716 173526 79744
rect 173590 79756 173618 79840
rect 173774 79824 173802 79908
rect 173710 79772 173716 79824
rect 173768 79784 173802 79824
rect 173768 79772 173774 79784
rect 173866 79756 173894 79988
rect 174418 79960 174446 80124
rect 178494 80112 178500 80124
rect 178552 80112 178558 80164
rect 177758 80044 177764 80096
rect 177816 80084 177822 80096
rect 181162 80084 181168 80096
rect 177816 80056 181168 80084
rect 177816 80044 177822 80056
rect 181162 80044 181168 80056
rect 181220 80044 181226 80096
rect 183526 80084 183554 80396
rect 238754 80084 238760 80096
rect 183526 80056 238760 80084
rect 238754 80044 238760 80056
rect 238812 80044 238818 80096
rect 177850 80016 177856 80028
rect 175614 79988 176286 80016
rect 173940 79908 173946 79960
rect 173998 79908 174004 79960
rect 174400 79908 174406 79960
rect 174458 79908 174464 79960
rect 174584 79908 174590 79960
rect 174642 79908 174648 79960
rect 174676 79908 174682 79960
rect 174734 79908 174740 79960
rect 174768 79908 174774 79960
rect 174826 79948 174832 79960
rect 174826 79920 175458 79948
rect 174826 79908 174832 79920
rect 173590 79716 173624 79756
rect 172848 79704 172854 79716
rect 173618 79704 173624 79716
rect 173676 79704 173682 79756
rect 173802 79704 173808 79756
rect 173860 79716 173894 79756
rect 173860 79704 173866 79716
rect 173958 79688 173986 79908
rect 174216 79840 174222 79892
rect 174274 79840 174280 79892
rect 174492 79840 174498 79892
rect 174550 79840 174556 79892
rect 171468 79648 171778 79676
rect 171468 79636 171474 79648
rect 173894 79636 173900 79688
rect 173952 79648 173986 79688
rect 174234 79676 174262 79840
rect 174354 79772 174360 79824
rect 174412 79812 174418 79824
rect 174510 79812 174538 79840
rect 174412 79784 174538 79812
rect 174412 79772 174418 79784
rect 174602 79756 174630 79908
rect 174694 79824 174722 79908
rect 174952 79840 174958 79892
rect 175010 79840 175016 79892
rect 175044 79840 175050 79892
rect 175102 79880 175108 79892
rect 175102 79840 175136 79880
rect 174694 79784 174728 79824
rect 174722 79772 174728 79784
rect 174780 79772 174786 79824
rect 174860 79772 174866 79824
rect 174918 79772 174924 79824
rect 174602 79716 174636 79756
rect 174630 79704 174636 79716
rect 174688 79704 174694 79756
rect 174878 79688 174906 79772
rect 174970 79756 174998 79840
rect 174970 79716 175004 79756
rect 174998 79704 175004 79716
rect 175056 79704 175062 79756
rect 175108 79688 175136 79840
rect 175430 79824 175458 79920
rect 175504 79908 175510 79960
rect 175562 79948 175568 79960
rect 175614 79948 175642 79988
rect 175964 79948 175970 79960
rect 175562 79920 175642 79948
rect 175562 79908 175568 79920
rect 175936 79908 175970 79948
rect 176022 79908 176028 79960
rect 176258 79948 176286 79988
rect 177086 79988 177856 80016
rect 177086 79960 177114 79988
rect 177850 79976 177856 79988
rect 177908 79976 177914 80028
rect 178586 80016 178592 80028
rect 178006 79988 178592 80016
rect 176258 79920 176470 79948
rect 175430 79784 175464 79824
rect 175458 79772 175464 79784
rect 175516 79772 175522 79824
rect 175596 79772 175602 79824
rect 175654 79772 175660 79824
rect 175688 79772 175694 79824
rect 175746 79812 175752 79824
rect 175746 79772 175780 79812
rect 175614 79688 175642 79772
rect 174538 79676 174544 79688
rect 174234 79648 174544 79676
rect 173952 79636 173958 79648
rect 174538 79636 174544 79648
rect 174596 79636 174602 79688
rect 174814 79636 174820 79688
rect 174872 79648 174906 79688
rect 174872 79636 174878 79648
rect 175090 79636 175096 79688
rect 175148 79636 175154 79688
rect 175614 79648 175648 79688
rect 175642 79636 175648 79648
rect 175700 79636 175706 79688
rect 171336 79580 174308 79608
rect 170456 79512 170628 79540
rect 171888 79512 173940 79540
rect 170456 79500 170462 79512
rect 171888 79472 171916 79512
rect 169444 79444 169984 79472
rect 171796 79444 171916 79472
rect 173912 79472 173940 79512
rect 174170 79472 174176 79484
rect 173912 79444 174176 79472
rect 169444 79432 169450 79444
rect 161624 79376 164556 79404
rect 161624 79364 161630 79376
rect 154758 79296 154764 79348
rect 154816 79336 154822 79348
rect 164418 79336 164424 79348
rect 154816 79308 164424 79336
rect 154816 79296 154822 79308
rect 164418 79296 164424 79308
rect 164476 79296 164482 79348
rect 164528 79336 164556 79376
rect 171686 79364 171692 79416
rect 171744 79404 171750 79416
rect 171796 79404 171824 79444
rect 174170 79432 174176 79444
rect 174228 79432 174234 79484
rect 174280 79472 174308 79580
rect 175274 79568 175280 79620
rect 175332 79608 175338 79620
rect 175752 79608 175780 79772
rect 175936 79688 175964 79908
rect 176148 79880 176154 79892
rect 176120 79840 176154 79880
rect 176206 79840 176212 79892
rect 176240 79840 176246 79892
rect 176298 79840 176304 79892
rect 176442 79880 176470 79920
rect 177068 79908 177074 79960
rect 177126 79908 177132 79960
rect 176442 79852 176562 79880
rect 175918 79636 175924 79688
rect 175976 79636 175982 79688
rect 176120 79620 176148 79840
rect 176258 79812 176286 79840
rect 176212 79784 176286 79812
rect 176212 79756 176240 79784
rect 176424 79772 176430 79824
rect 176482 79772 176488 79824
rect 176194 79704 176200 79756
rect 176252 79704 176258 79756
rect 176286 79704 176292 79756
rect 176344 79744 176350 79756
rect 176442 79744 176470 79772
rect 176344 79716 176470 79744
rect 176344 79704 176350 79716
rect 176378 79636 176384 79688
rect 176436 79676 176442 79688
rect 176534 79676 176562 79852
rect 176792 79840 176798 79892
rect 176850 79880 176856 79892
rect 177850 79880 177856 79892
rect 176850 79852 177856 79880
rect 176850 79840 176856 79852
rect 177850 79840 177856 79852
rect 177908 79840 177914 79892
rect 176700 79772 176706 79824
rect 176758 79772 176764 79824
rect 177574 79772 177580 79824
rect 177632 79812 177638 79824
rect 178006 79812 178034 79988
rect 178586 79976 178592 79988
rect 178644 79976 178650 80028
rect 177632 79784 178034 79812
rect 177632 79772 177638 79784
rect 176436 79648 176562 79676
rect 176718 79676 176746 79772
rect 178218 79704 178224 79756
rect 178276 79744 178282 79756
rect 191282 79744 191288 79756
rect 178276 79716 191288 79744
rect 178276 79704 178282 79716
rect 191282 79704 191288 79716
rect 191340 79704 191346 79756
rect 176718 79648 176792 79676
rect 176436 79636 176442 79648
rect 175332 79580 175780 79608
rect 175332 79568 175338 79580
rect 176102 79568 176108 79620
rect 176160 79568 176166 79620
rect 176764 79552 176792 79648
rect 178126 79636 178132 79688
rect 178184 79676 178190 79688
rect 189810 79676 189816 79688
rect 178184 79648 189816 79676
rect 178184 79636 178190 79648
rect 189810 79636 189816 79648
rect 189868 79636 189874 79688
rect 177482 79568 177488 79620
rect 177540 79608 177546 79620
rect 190730 79608 190736 79620
rect 177540 79580 190736 79608
rect 177540 79568 177546 79580
rect 190730 79568 190736 79580
rect 190788 79608 190794 79620
rect 190788 79580 200114 79608
rect 190788 79568 190794 79580
rect 175366 79500 175372 79552
rect 175424 79540 175430 79552
rect 175826 79540 175832 79552
rect 175424 79512 175832 79540
rect 175424 79500 175430 79512
rect 175826 79500 175832 79512
rect 175884 79500 175890 79552
rect 176746 79500 176752 79552
rect 176804 79500 176810 79552
rect 178770 79540 178776 79552
rect 176856 79512 178776 79540
rect 176856 79472 176884 79512
rect 178770 79500 178776 79512
rect 178828 79500 178834 79552
rect 174280 79444 176884 79472
rect 178034 79432 178040 79484
rect 178092 79472 178098 79484
rect 194042 79472 194048 79484
rect 178092 79444 194048 79472
rect 178092 79432 178098 79444
rect 194042 79432 194048 79444
rect 194100 79432 194106 79484
rect 200086 79404 200114 79580
rect 306374 79404 306380 79416
rect 171744 79376 171824 79404
rect 171888 79376 179414 79404
rect 200086 79376 306380 79404
rect 171744 79364 171750 79376
rect 171888 79336 171916 79376
rect 164528 79308 171916 79336
rect 171980 79308 173710 79336
rect 163958 79268 163964 79280
rect 154546 79240 163964 79268
rect 163958 79228 163964 79240
rect 164016 79228 164022 79280
rect 165706 79228 165712 79280
rect 165764 79268 165770 79280
rect 165890 79268 165896 79280
rect 165764 79240 165896 79268
rect 165764 79228 165770 79240
rect 165890 79228 165896 79240
rect 165948 79268 165954 79280
rect 171980 79268 172008 79308
rect 173682 79268 173710 79308
rect 174354 79296 174360 79348
rect 174412 79336 174418 79348
rect 177758 79336 177764 79348
rect 174412 79308 177764 79336
rect 174412 79296 174418 79308
rect 177758 79296 177764 79308
rect 177816 79296 177822 79348
rect 179386 79336 179414 79376
rect 306374 79364 306380 79376
rect 306432 79364 306438 79416
rect 189902 79336 189908 79348
rect 179386 79308 189908 79336
rect 189902 79296 189908 79308
rect 189960 79296 189966 79348
rect 324314 79336 324320 79348
rect 200086 79308 324320 79336
rect 193858 79268 193864 79280
rect 165948 79240 172008 79268
rect 173498 79240 173618 79268
rect 173682 79240 193864 79268
rect 165948 79228 165954 79240
rect 143040 79172 153194 79200
rect 143040 79160 143046 79172
rect 167362 79160 167368 79212
rect 167420 79200 167426 79212
rect 173498 79200 173526 79240
rect 167420 79172 173526 79200
rect 173590 79200 173618 79240
rect 193858 79228 193864 79240
rect 193916 79228 193922 79280
rect 196802 79200 196808 79212
rect 173590 79172 196808 79200
rect 167420 79160 167426 79172
rect 196802 79160 196808 79172
rect 196860 79160 196866 79212
rect 147398 79132 147404 79144
rect 120684 79104 141924 79132
rect 141988 79104 147404 79132
rect 120684 79092 120690 79104
rect 119246 79024 119252 79076
rect 119304 79064 119310 79076
rect 141988 79064 142016 79104
rect 147398 79092 147404 79104
rect 147456 79092 147462 79144
rect 160646 79092 160652 79144
rect 160704 79132 160710 79144
rect 192938 79132 192944 79144
rect 160704 79104 173296 79132
rect 160704 79092 160710 79104
rect 147214 79064 147220 79076
rect 119304 79036 142016 79064
rect 142080 79036 147220 79064
rect 119304 79024 119310 79036
rect 118050 78956 118056 79008
rect 118108 78996 118114 79008
rect 142080 78996 142108 79036
rect 147214 79024 147220 79036
rect 147272 79024 147278 79076
rect 157610 79024 157616 79076
rect 157668 79064 157674 79076
rect 173158 79064 173164 79076
rect 157668 79036 173164 79064
rect 157668 79024 157674 79036
rect 173158 79024 173164 79036
rect 173216 79024 173222 79076
rect 173268 79064 173296 79104
rect 173636 79104 192944 79132
rect 173636 79064 173664 79104
rect 192938 79092 192944 79104
rect 192996 79092 193002 79144
rect 173268 79036 173664 79064
rect 173802 79024 173808 79076
rect 173860 79064 173866 79076
rect 192018 79064 192024 79076
rect 173860 79036 192024 79064
rect 173860 79024 173866 79036
rect 192018 79024 192024 79036
rect 192076 79064 192082 79076
rect 200086 79064 200114 79308
rect 324314 79296 324320 79308
rect 324372 79296 324378 79348
rect 192076 79036 200114 79064
rect 192076 79024 192082 79036
rect 118108 78968 142108 78996
rect 118108 78956 118114 78968
rect 142154 78956 142160 79008
rect 142212 78996 142218 79008
rect 147858 78996 147864 79008
rect 142212 78968 147864 78996
rect 142212 78956 142218 78968
rect 147858 78956 147864 78968
rect 147916 78956 147922 79008
rect 168098 78956 168104 79008
rect 168156 78996 168162 79008
rect 168282 78996 168288 79008
rect 168156 78968 168288 78996
rect 168156 78956 168162 78968
rect 168282 78956 168288 78968
rect 168340 78996 168346 79008
rect 201862 78996 201868 79008
rect 168340 78968 201868 78996
rect 168340 78956 168346 78968
rect 201862 78956 201868 78968
rect 201920 78956 201926 79008
rect 117590 78888 117596 78940
rect 117648 78928 117654 78940
rect 140498 78928 140504 78940
rect 117648 78900 140504 78928
rect 117648 78888 117654 78900
rect 140498 78888 140504 78900
rect 140556 78888 140562 78940
rect 141326 78888 141332 78940
rect 141384 78928 141390 78940
rect 145374 78928 145380 78940
rect 141384 78900 145380 78928
rect 141384 78888 141390 78900
rect 145374 78888 145380 78900
rect 145432 78888 145438 78940
rect 148686 78888 148692 78940
rect 148744 78928 148750 78940
rect 148744 78900 154712 78928
rect 148744 78888 148750 78900
rect 117866 78820 117872 78872
rect 117924 78860 117930 78872
rect 154684 78860 154712 78900
rect 157610 78888 157616 78940
rect 157668 78928 157674 78940
rect 157794 78928 157800 78940
rect 157668 78900 157800 78928
rect 157668 78888 157674 78900
rect 157794 78888 157800 78900
rect 157852 78888 157858 78940
rect 163958 78888 163964 78940
rect 164016 78928 164022 78940
rect 169018 78928 169024 78940
rect 164016 78900 169024 78928
rect 164016 78888 164022 78900
rect 169018 78888 169024 78900
rect 169076 78888 169082 78940
rect 169202 78888 169208 78940
rect 169260 78928 169266 78940
rect 170858 78928 170864 78940
rect 169260 78900 170864 78928
rect 169260 78888 169266 78900
rect 170858 78888 170864 78900
rect 170916 78888 170922 78940
rect 171502 78888 171508 78940
rect 171560 78928 171566 78940
rect 172146 78928 172152 78940
rect 171560 78900 172152 78928
rect 171560 78888 171566 78900
rect 172146 78888 172152 78900
rect 172204 78888 172210 78940
rect 172606 78888 172612 78940
rect 172664 78928 172670 78940
rect 181070 78928 181076 78940
rect 172664 78900 181076 78928
rect 172664 78888 172670 78900
rect 181070 78888 181076 78900
rect 181128 78928 181134 78940
rect 288434 78928 288440 78940
rect 181128 78900 288440 78928
rect 181128 78888 181134 78900
rect 288434 78888 288440 78900
rect 288492 78888 288498 78940
rect 180886 78860 180892 78872
rect 117924 78832 140176 78860
rect 117924 78820 117930 78832
rect 130102 78752 130108 78804
rect 130160 78792 130166 78804
rect 140038 78792 140044 78804
rect 130160 78764 140044 78792
rect 130160 78752 130166 78764
rect 140038 78752 140044 78764
rect 140096 78752 140102 78804
rect 140148 78792 140176 78832
rect 142310 78832 149100 78860
rect 154684 78832 180892 78860
rect 142310 78792 142338 78832
rect 149072 78804 149100 78832
rect 180886 78820 180892 78832
rect 180944 78820 180950 78872
rect 186314 78820 186320 78872
rect 186372 78860 186378 78872
rect 186958 78860 186964 78872
rect 186372 78832 186964 78860
rect 186372 78820 186378 78832
rect 186958 78820 186964 78832
rect 187016 78860 187022 78872
rect 480254 78860 480260 78872
rect 187016 78832 480260 78860
rect 187016 78820 187022 78832
rect 480254 78820 480260 78832
rect 480312 78820 480318 78872
rect 140148 78764 142338 78792
rect 149054 78752 149060 78804
rect 149112 78792 149118 78804
rect 150066 78792 150072 78804
rect 149112 78764 150072 78792
rect 149112 78752 149118 78764
rect 150066 78752 150072 78764
rect 150124 78752 150130 78804
rect 151998 78752 152004 78804
rect 152056 78792 152062 78804
rect 152182 78792 152188 78804
rect 152056 78764 152188 78792
rect 152056 78752 152062 78764
rect 152182 78752 152188 78764
rect 152240 78752 152246 78804
rect 170306 78752 170312 78804
rect 170364 78792 170370 78804
rect 172606 78792 172612 78804
rect 170364 78764 172612 78792
rect 170364 78752 170370 78764
rect 172606 78752 172612 78764
rect 172664 78752 172670 78804
rect 173158 78752 173164 78804
rect 173216 78792 173222 78804
rect 173802 78792 173808 78804
rect 173216 78764 173808 78792
rect 173216 78752 173222 78764
rect 173802 78752 173808 78764
rect 173860 78752 173866 78804
rect 173986 78752 173992 78804
rect 174044 78792 174050 78804
rect 178218 78792 178224 78804
rect 174044 78764 178224 78792
rect 174044 78752 174050 78764
rect 178218 78752 178224 78764
rect 178276 78752 178282 78804
rect 186406 78752 186412 78804
rect 186464 78792 186470 78804
rect 187050 78792 187056 78804
rect 186464 78764 187056 78792
rect 186464 78752 186470 78764
rect 187050 78752 187056 78764
rect 187108 78792 187114 78804
rect 483014 78792 483020 78804
rect 187108 78764 483020 78792
rect 187108 78752 187114 78764
rect 483014 78752 483020 78764
rect 483072 78752 483078 78804
rect 131850 78684 131856 78736
rect 131908 78724 131914 78736
rect 137554 78724 137560 78736
rect 131908 78696 137560 78724
rect 131908 78684 131914 78696
rect 137554 78684 137560 78696
rect 137612 78684 137618 78736
rect 140958 78684 140964 78736
rect 141016 78724 141022 78736
rect 141326 78724 141332 78736
rect 141016 78696 141332 78724
rect 141016 78684 141022 78696
rect 141326 78684 141332 78696
rect 141384 78684 141390 78736
rect 146846 78684 146852 78736
rect 146904 78724 146910 78736
rect 179506 78724 179512 78736
rect 146904 78696 179512 78724
rect 146904 78684 146910 78696
rect 179506 78684 179512 78696
rect 179564 78684 179570 78736
rect 187694 78684 187700 78736
rect 187752 78724 187758 78736
rect 188338 78724 188344 78736
rect 187752 78696 188344 78724
rect 187752 78684 187758 78696
rect 188338 78684 188344 78696
rect 188396 78724 188402 78736
rect 500954 78724 500960 78736
rect 188396 78696 500960 78724
rect 188396 78684 188402 78696
rect 500954 78684 500960 78696
rect 501012 78684 501018 78736
rect 120074 78616 120080 78668
rect 120132 78656 120138 78668
rect 121362 78656 121368 78668
rect 120132 78628 121368 78656
rect 120132 78616 120138 78628
rect 121362 78616 121368 78628
rect 121420 78656 121426 78668
rect 132034 78656 132040 78668
rect 121420 78628 132040 78656
rect 121420 78616 121426 78628
rect 132034 78616 132040 78628
rect 132092 78616 132098 78668
rect 133690 78616 133696 78668
rect 133748 78656 133754 78668
rect 133874 78656 133880 78668
rect 133748 78628 133880 78656
rect 133748 78616 133754 78628
rect 133874 78616 133880 78628
rect 133932 78616 133938 78668
rect 138382 78616 138388 78668
rect 138440 78656 138446 78668
rect 138566 78656 138572 78668
rect 138440 78628 138572 78656
rect 138440 78616 138446 78628
rect 138566 78616 138572 78628
rect 138624 78616 138630 78668
rect 138842 78616 138848 78668
rect 138900 78656 138906 78668
rect 139118 78656 139124 78668
rect 138900 78628 139124 78656
rect 138900 78616 138906 78628
rect 139118 78616 139124 78628
rect 139176 78616 139182 78668
rect 140498 78616 140504 78668
rect 140556 78656 140562 78668
rect 146294 78656 146300 78668
rect 140556 78628 146300 78656
rect 140556 78616 140562 78628
rect 146294 78616 146300 78628
rect 146352 78656 146358 78668
rect 148962 78656 148968 78668
rect 146352 78628 148968 78656
rect 146352 78616 146358 78628
rect 148962 78616 148968 78628
rect 149020 78616 149026 78668
rect 151998 78616 152004 78668
rect 152056 78656 152062 78668
rect 152366 78656 152372 78668
rect 152056 78628 152372 78656
rect 152056 78616 152062 78628
rect 152366 78616 152372 78628
rect 152424 78616 152430 78668
rect 153286 78616 153292 78668
rect 153344 78656 153350 78668
rect 154114 78656 154120 78668
rect 153344 78628 154120 78656
rect 153344 78616 153350 78628
rect 154114 78616 154120 78628
rect 154172 78616 154178 78668
rect 165798 78616 165804 78668
rect 165856 78656 165862 78668
rect 196250 78656 196256 78668
rect 165856 78628 196256 78656
rect 165856 78616 165862 78628
rect 196250 78616 196256 78628
rect 196308 78656 196314 78668
rect 196618 78656 196624 78668
rect 196308 78628 196624 78656
rect 196308 78616 196314 78628
rect 196618 78616 196624 78628
rect 196676 78616 196682 78668
rect 102134 78548 102140 78600
rect 102192 78588 102198 78600
rect 102778 78588 102784 78600
rect 102192 78560 102784 78588
rect 102192 78548 102198 78560
rect 102778 78548 102784 78560
rect 102836 78588 102842 78600
rect 134058 78588 134064 78600
rect 102836 78560 134064 78588
rect 102836 78548 102842 78560
rect 134058 78548 134064 78560
rect 134116 78548 134122 78600
rect 137554 78548 137560 78600
rect 137612 78588 137618 78600
rect 143350 78588 143356 78600
rect 137612 78560 143356 78588
rect 137612 78548 137618 78560
rect 143350 78548 143356 78560
rect 143408 78548 143414 78600
rect 147214 78548 147220 78600
rect 147272 78588 147278 78600
rect 150526 78588 150532 78600
rect 147272 78560 150532 78588
rect 147272 78548 147278 78560
rect 150526 78548 150532 78560
rect 150584 78548 150590 78600
rect 164418 78548 164424 78600
rect 164476 78588 164482 78600
rect 164476 78560 168972 78588
rect 164476 78548 164482 78560
rect 130838 78480 130844 78532
rect 130896 78520 130902 78532
rect 133874 78520 133880 78532
rect 130896 78492 133880 78520
rect 130896 78480 130902 78492
rect 133874 78480 133880 78492
rect 133932 78480 133938 78532
rect 142614 78520 142620 78532
rect 135226 78492 142620 78520
rect 104066 78412 104072 78464
rect 104124 78452 104130 78464
rect 130470 78452 130476 78464
rect 104124 78424 130476 78452
rect 104124 78412 104130 78424
rect 130470 78412 130476 78424
rect 130528 78412 130534 78464
rect 132586 78344 132592 78396
rect 132644 78384 132650 78396
rect 135226 78384 135254 78492
rect 142614 78480 142620 78492
rect 142672 78480 142678 78532
rect 142982 78480 142988 78532
rect 143040 78480 143046 78532
rect 168944 78520 168972 78560
rect 169662 78548 169668 78600
rect 169720 78588 169726 78600
rect 169720 78560 173894 78588
rect 169720 78548 169726 78560
rect 170306 78520 170312 78532
rect 168944 78492 170312 78520
rect 170306 78480 170312 78492
rect 170364 78480 170370 78532
rect 171870 78480 171876 78532
rect 171928 78520 171934 78532
rect 172238 78520 172244 78532
rect 171928 78492 172244 78520
rect 171928 78480 171934 78492
rect 172238 78480 172244 78492
rect 172296 78480 172302 78532
rect 173866 78520 173894 78560
rect 181438 78548 181444 78600
rect 181496 78588 181502 78600
rect 192846 78588 192852 78600
rect 181496 78560 192852 78588
rect 181496 78548 181502 78560
rect 192846 78548 192852 78560
rect 192904 78548 192910 78600
rect 186314 78520 186320 78532
rect 173866 78492 186320 78520
rect 186314 78480 186320 78492
rect 186372 78480 186378 78532
rect 137094 78412 137100 78464
rect 137152 78452 137158 78464
rect 142062 78452 142068 78464
rect 137152 78424 142068 78452
rect 137152 78412 137158 78424
rect 142062 78412 142068 78424
rect 142120 78412 142126 78464
rect 143000 78452 143028 78480
rect 142632 78424 143028 78452
rect 142632 78396 142660 78424
rect 153746 78412 153752 78464
rect 153804 78452 153810 78464
rect 154482 78452 154488 78464
rect 153804 78424 154488 78452
rect 153804 78412 153810 78424
rect 154482 78412 154488 78424
rect 154540 78412 154546 78464
rect 158806 78412 158812 78464
rect 158864 78452 158870 78464
rect 163406 78452 163412 78464
rect 158864 78424 163412 78452
rect 158864 78412 158870 78424
rect 163406 78412 163412 78424
rect 163464 78412 163470 78464
rect 170030 78412 170036 78464
rect 170088 78452 170094 78464
rect 186406 78452 186412 78464
rect 170088 78424 186412 78452
rect 170088 78412 170094 78424
rect 186406 78412 186412 78424
rect 186464 78412 186470 78464
rect 132644 78356 135254 78384
rect 132644 78344 132650 78356
rect 139118 78344 139124 78396
rect 139176 78384 139182 78396
rect 139302 78384 139308 78396
rect 139176 78356 139308 78384
rect 139176 78344 139182 78356
rect 139302 78344 139308 78356
rect 139360 78344 139366 78396
rect 140958 78344 140964 78396
rect 141016 78384 141022 78396
rect 141418 78384 141424 78396
rect 141016 78356 141424 78384
rect 141016 78344 141022 78356
rect 141418 78344 141424 78356
rect 141476 78344 141482 78396
rect 142614 78344 142620 78396
rect 142672 78344 142678 78396
rect 142982 78344 142988 78396
rect 143040 78384 143046 78396
rect 143534 78384 143540 78396
rect 143040 78356 143540 78384
rect 143040 78344 143046 78356
rect 143534 78344 143540 78356
rect 143592 78344 143598 78396
rect 163222 78344 163228 78396
rect 163280 78384 163286 78396
rect 164142 78384 164148 78396
rect 163280 78356 164148 78384
rect 163280 78344 163286 78356
rect 164142 78344 164148 78356
rect 164200 78344 164206 78396
rect 165890 78344 165896 78396
rect 165948 78384 165954 78396
rect 166166 78384 166172 78396
rect 165948 78356 166172 78384
rect 165948 78344 165954 78356
rect 166166 78344 166172 78356
rect 166224 78344 166230 78396
rect 166994 78344 167000 78396
rect 167052 78384 167058 78396
rect 183094 78384 183100 78396
rect 167052 78356 183100 78384
rect 167052 78344 167058 78356
rect 183094 78344 183100 78356
rect 183152 78344 183158 78396
rect 205818 78344 205824 78396
rect 205876 78384 205882 78396
rect 206186 78384 206192 78396
rect 205876 78356 206192 78384
rect 205876 78344 205882 78356
rect 206186 78344 206192 78356
rect 206244 78344 206250 78396
rect 57974 78276 57980 78328
rect 58032 78316 58038 78328
rect 107286 78316 107292 78328
rect 58032 78288 107292 78316
rect 58032 78276 58038 78288
rect 107286 78276 107292 78288
rect 107344 78276 107350 78328
rect 122190 78276 122196 78328
rect 122248 78316 122254 78328
rect 148502 78316 148508 78328
rect 122248 78288 148508 78316
rect 122248 78276 122254 78288
rect 148502 78276 148508 78288
rect 148560 78276 148566 78328
rect 167454 78276 167460 78328
rect 167512 78316 167518 78328
rect 253198 78316 253204 78328
rect 167512 78288 253204 78316
rect 167512 78276 167518 78288
rect 253198 78276 253204 78288
rect 253256 78276 253262 78328
rect 46934 78208 46940 78260
rect 46992 78248 46998 78260
rect 107194 78248 107200 78260
rect 46992 78220 107200 78248
rect 46992 78208 46998 78220
rect 107194 78208 107200 78220
rect 107252 78208 107258 78260
rect 123386 78208 123392 78260
rect 123444 78248 123450 78260
rect 123444 78220 138198 78248
rect 123444 78208 123450 78220
rect 20714 78140 20720 78192
rect 20772 78180 20778 78192
rect 102134 78180 102140 78192
rect 20772 78152 102140 78180
rect 20772 78140 20778 78152
rect 102134 78140 102140 78152
rect 102192 78140 102198 78192
rect 130194 78180 130200 78192
rect 113146 78152 130200 78180
rect 6914 78072 6920 78124
rect 6972 78112 6978 78124
rect 107102 78112 107108 78124
rect 6972 78084 107108 78112
rect 6972 78072 6978 78084
rect 107102 78072 107108 78084
rect 107160 78112 107166 78124
rect 107378 78112 107384 78124
rect 107160 78084 107384 78112
rect 107160 78072 107166 78084
rect 107378 78072 107384 78084
rect 107436 78072 107442 78124
rect 2774 78004 2780 78056
rect 2832 78044 2838 78056
rect 104066 78044 104072 78056
rect 2832 78016 104072 78044
rect 2832 78004 2838 78016
rect 104066 78004 104072 78016
rect 104124 78004 104130 78056
rect 2866 77936 2872 77988
rect 2924 77976 2930 77988
rect 108574 77976 108580 77988
rect 2924 77948 108580 77976
rect 2924 77936 2930 77948
rect 108574 77936 108580 77948
rect 108632 77976 108638 77988
rect 113146 77976 113174 78152
rect 130194 78140 130200 78152
rect 130252 78140 130258 78192
rect 133874 78140 133880 78192
rect 133932 78180 133938 78192
rect 137554 78180 137560 78192
rect 133932 78152 137560 78180
rect 133932 78140 133938 78152
rect 137554 78140 137560 78152
rect 137612 78140 137618 78192
rect 138170 78180 138198 78220
rect 138290 78208 138296 78260
rect 138348 78248 138354 78260
rect 144086 78248 144092 78260
rect 138348 78220 144092 78248
rect 138348 78208 138354 78220
rect 144086 78208 144092 78220
rect 144144 78208 144150 78260
rect 150618 78208 150624 78260
rect 150676 78248 150682 78260
rect 151170 78248 151176 78260
rect 150676 78220 151176 78248
rect 150676 78208 150682 78220
rect 151170 78208 151176 78220
rect 151228 78208 151234 78260
rect 160922 78208 160928 78260
rect 160980 78248 160986 78260
rect 166166 78248 166172 78260
rect 160980 78220 166172 78248
rect 160980 78208 160986 78220
rect 166166 78208 166172 78220
rect 166224 78208 166230 78260
rect 169846 78208 169852 78260
rect 169904 78208 169910 78260
rect 170858 78208 170864 78260
rect 170916 78248 170922 78260
rect 337378 78248 337384 78260
rect 170916 78220 337384 78248
rect 170916 78208 170922 78220
rect 337378 78208 337384 78220
rect 337436 78208 337442 78260
rect 148318 78180 148324 78192
rect 138170 78152 148324 78180
rect 148318 78140 148324 78152
rect 148376 78140 148382 78192
rect 152550 78140 152556 78192
rect 152608 78180 152614 78192
rect 153010 78180 153016 78192
rect 152608 78152 153016 78180
rect 152608 78140 152614 78152
rect 153010 78140 153016 78152
rect 153068 78140 153074 78192
rect 161474 78140 161480 78192
rect 161532 78180 161538 78192
rect 162026 78180 162032 78192
rect 161532 78152 162032 78180
rect 161532 78140 161538 78152
rect 162026 78140 162032 78152
rect 162084 78140 162090 78192
rect 169864 78180 169892 78208
rect 400858 78180 400864 78192
rect 169864 78152 400864 78180
rect 400858 78140 400864 78152
rect 400916 78140 400922 78192
rect 123018 78072 123024 78124
rect 123076 78112 123082 78124
rect 143442 78112 143448 78124
rect 123076 78084 143448 78112
rect 123076 78072 123082 78084
rect 143442 78072 143448 78084
rect 143500 78072 143506 78124
rect 149698 78072 149704 78124
rect 149756 78112 149762 78124
rect 183646 78112 183652 78124
rect 149756 78084 183652 78112
rect 149756 78072 149762 78084
rect 183646 78072 183652 78084
rect 183704 78072 183710 78124
rect 196250 78072 196256 78124
rect 196308 78112 196314 78124
rect 429194 78112 429200 78124
rect 196308 78084 429200 78112
rect 196308 78072 196314 78084
rect 429194 78072 429200 78084
rect 429252 78072 429258 78124
rect 113634 78004 113640 78056
rect 113692 78044 113698 78056
rect 129826 78044 129832 78056
rect 113692 78016 129832 78044
rect 113692 78004 113698 78016
rect 129826 78004 129832 78016
rect 129884 78044 129890 78056
rect 131850 78044 131856 78056
rect 129884 78016 131856 78044
rect 129884 78004 129890 78016
rect 131850 78004 131856 78016
rect 131908 78004 131914 78056
rect 173986 78044 173992 78056
rect 162872 78016 173992 78044
rect 108632 77948 113174 77976
rect 108632 77936 108638 77948
rect 132494 77936 132500 77988
rect 132552 77976 132558 77988
rect 137094 77976 137100 77988
rect 132552 77948 137100 77976
rect 132552 77936 132558 77948
rect 137094 77936 137100 77948
rect 137152 77936 137158 77988
rect 153194 77936 153200 77988
rect 153252 77976 153258 77988
rect 153654 77976 153660 77988
rect 153252 77948 153660 77976
rect 153252 77936 153258 77948
rect 153654 77936 153660 77948
rect 153712 77936 153718 77988
rect 156414 77936 156420 77988
rect 156472 77976 156478 77988
rect 161474 77976 161480 77988
rect 156472 77948 161480 77976
rect 156472 77936 156478 77948
rect 161474 77936 161480 77948
rect 161532 77936 161538 77988
rect 131022 77868 131028 77920
rect 131080 77908 131086 77920
rect 142522 77908 142528 77920
rect 131080 77880 142528 77908
rect 131080 77868 131086 77880
rect 142522 77868 142528 77880
rect 142580 77868 142586 77920
rect 148410 77868 148416 77920
rect 148468 77908 148474 77920
rect 148778 77908 148784 77920
rect 148468 77880 148784 77908
rect 148468 77868 148474 77880
rect 148778 77868 148784 77880
rect 148836 77868 148842 77920
rect 107378 77800 107384 77852
rect 107436 77840 107442 77852
rect 129458 77840 129464 77852
rect 107436 77812 129464 77840
rect 107436 77800 107442 77812
rect 129458 77800 129464 77812
rect 129516 77800 129522 77852
rect 129550 77800 129556 77852
rect 129608 77840 129614 77852
rect 134426 77840 134432 77852
rect 129608 77812 134432 77840
rect 129608 77800 129614 77812
rect 134426 77800 134432 77812
rect 134484 77800 134490 77852
rect 150434 77840 150440 77852
rect 137986 77812 150440 77840
rect 131942 77732 131948 77784
rect 132000 77772 132006 77784
rect 137986 77772 138014 77812
rect 150434 77800 150440 77812
rect 150492 77840 150498 77852
rect 151446 77840 151452 77852
rect 150492 77812 151452 77840
rect 150492 77800 150498 77812
rect 151446 77800 151452 77812
rect 151504 77800 151510 77852
rect 157426 77800 157432 77852
rect 157484 77840 157490 77852
rect 157794 77840 157800 77852
rect 157484 77812 157800 77840
rect 157484 77800 157490 77812
rect 157794 77800 157800 77812
rect 157852 77800 157858 77852
rect 132000 77744 138014 77772
rect 132000 77732 132006 77744
rect 159358 77732 159364 77784
rect 159416 77772 159422 77784
rect 162872 77772 162900 78016
rect 173986 78004 173992 78016
rect 174044 78004 174050 78056
rect 174170 78004 174176 78056
rect 174228 78044 174234 78056
rect 178954 78044 178960 78056
rect 174228 78016 178960 78044
rect 174228 78004 174234 78016
rect 178954 78004 178960 78016
rect 179012 78004 179018 78056
rect 180794 78004 180800 78056
rect 180852 78044 180858 78056
rect 415486 78044 415492 78056
rect 180852 78016 415492 78044
rect 180852 78004 180858 78016
rect 415486 78004 415492 78016
rect 415544 78004 415550 78056
rect 169478 77936 169484 77988
rect 169536 77976 169542 77988
rect 169754 77976 169760 77988
rect 169536 77948 169760 77976
rect 169536 77936 169542 77948
rect 169754 77936 169760 77948
rect 169812 77936 169818 77988
rect 177390 77936 177396 77988
rect 177448 77976 177454 77988
rect 177850 77976 177856 77988
rect 177448 77948 177856 77976
rect 177448 77936 177454 77948
rect 177850 77936 177856 77948
rect 177908 77936 177914 77988
rect 422294 77976 422300 77988
rect 179386 77948 422300 77976
rect 162946 77868 162952 77920
rect 163004 77908 163010 77920
rect 177206 77908 177212 77920
rect 163004 77880 177212 77908
rect 163004 77868 163010 77880
rect 177206 77868 177212 77880
rect 177264 77868 177270 77920
rect 163498 77800 163504 77852
rect 163556 77840 163562 77852
rect 178770 77840 178776 77852
rect 163556 77812 178776 77840
rect 163556 77800 163562 77812
rect 178770 77800 178776 77812
rect 178828 77800 178834 77852
rect 159416 77744 162900 77772
rect 159416 77732 159422 77744
rect 165246 77732 165252 77784
rect 165304 77772 165310 77784
rect 179386 77772 179414 77948
rect 422294 77936 422300 77948
rect 422352 77936 422358 77988
rect 181530 77868 181536 77920
rect 181588 77908 181594 77920
rect 194134 77908 194140 77920
rect 181588 77880 194140 77908
rect 181588 77868 181594 77880
rect 194134 77868 194140 77880
rect 194192 77868 194198 77920
rect 165304 77744 179414 77772
rect 165304 77732 165310 77744
rect 107286 77664 107292 77716
rect 107344 77704 107350 77716
rect 136818 77704 136824 77716
rect 107344 77676 136824 77704
rect 107344 77664 107350 77676
rect 136818 77664 136824 77676
rect 136876 77664 136882 77716
rect 137094 77664 137100 77716
rect 137152 77704 137158 77716
rect 142338 77704 142344 77716
rect 137152 77676 142344 77704
rect 137152 77664 137158 77676
rect 142338 77664 142344 77676
rect 142396 77664 142402 77716
rect 169846 77664 169852 77716
rect 169904 77704 169910 77716
rect 171134 77704 171140 77716
rect 169904 77676 171140 77704
rect 169904 77664 169910 77676
rect 171134 77664 171140 77676
rect 171192 77704 171198 77716
rect 187510 77704 187516 77716
rect 171192 77676 187516 77704
rect 171192 77664 171198 77676
rect 187510 77664 187516 77676
rect 187568 77664 187574 77716
rect 131206 77596 131212 77648
rect 131264 77636 131270 77648
rect 132310 77636 132316 77648
rect 131264 77608 132316 77636
rect 131264 77596 131270 77608
rect 132310 77596 132316 77608
rect 132368 77636 132374 77648
rect 139854 77636 139860 77648
rect 132368 77608 139860 77636
rect 132368 77596 132374 77608
rect 139854 77596 139860 77608
rect 139912 77596 139918 77648
rect 156138 77596 156144 77648
rect 156196 77636 156202 77648
rect 162210 77636 162216 77648
rect 156196 77608 162216 77636
rect 156196 77596 156202 77608
rect 162210 77596 162216 77608
rect 162268 77596 162274 77648
rect 131758 77528 131764 77580
rect 131816 77568 131822 77580
rect 142246 77568 142252 77580
rect 131816 77540 142252 77568
rect 131816 77528 131822 77540
rect 142246 77528 142252 77540
rect 142304 77528 142310 77580
rect 164602 77528 164608 77580
rect 164660 77568 164666 77580
rect 180794 77568 180800 77580
rect 164660 77540 180800 77568
rect 164660 77528 164666 77540
rect 180794 77528 180800 77540
rect 180852 77528 180858 77580
rect 107194 77460 107200 77512
rect 107252 77500 107258 77512
rect 136082 77500 136088 77512
rect 107252 77472 136088 77500
rect 107252 77460 107258 77472
rect 136082 77460 136088 77472
rect 136140 77460 136146 77512
rect 137002 77460 137008 77512
rect 137060 77500 137066 77512
rect 137370 77500 137376 77512
rect 137060 77472 137376 77500
rect 137060 77460 137066 77472
rect 137370 77460 137376 77472
rect 137428 77460 137434 77512
rect 164050 77460 164056 77512
rect 164108 77500 164114 77512
rect 178862 77500 178868 77512
rect 164108 77472 178868 77500
rect 164108 77460 164114 77472
rect 178862 77460 178868 77472
rect 178920 77460 178926 77512
rect 134058 77392 134064 77444
rect 134116 77432 134122 77444
rect 137554 77432 137560 77444
rect 134116 77404 137560 77432
rect 134116 77392 134122 77404
rect 137554 77392 137560 77404
rect 137612 77392 137618 77444
rect 138106 77392 138112 77444
rect 138164 77432 138170 77444
rect 146018 77432 146024 77444
rect 138164 77404 146024 77432
rect 138164 77392 138170 77404
rect 146018 77392 146024 77404
rect 146076 77392 146082 77444
rect 158346 77392 158352 77444
rect 158404 77432 158410 77444
rect 163498 77432 163504 77444
rect 158404 77404 163504 77432
rect 158404 77392 158410 77404
rect 163498 77392 163504 77404
rect 163556 77392 163562 77444
rect 164694 77392 164700 77444
rect 164752 77432 164758 77444
rect 165062 77432 165068 77444
rect 164752 77404 165068 77432
rect 164752 77392 164758 77404
rect 165062 77392 165068 77404
rect 165120 77432 165126 77444
rect 181438 77432 181444 77444
rect 165120 77404 181444 77432
rect 165120 77392 165126 77404
rect 181438 77392 181444 77404
rect 181496 77392 181502 77444
rect 130194 77324 130200 77376
rect 130252 77364 130258 77376
rect 133598 77364 133604 77376
rect 130252 77336 133604 77364
rect 130252 77324 130258 77336
rect 133598 77324 133604 77336
rect 133656 77324 133662 77376
rect 154850 77324 154856 77376
rect 154908 77364 154914 77376
rect 158622 77364 158628 77376
rect 154908 77336 158628 77364
rect 154908 77324 154914 77336
rect 158622 77324 158628 77336
rect 158680 77324 158686 77376
rect 160738 77324 160744 77376
rect 160796 77364 160802 77376
rect 161382 77364 161388 77376
rect 160796 77336 161388 77364
rect 160796 77324 160802 77336
rect 161382 77324 161388 77336
rect 161440 77324 161446 77376
rect 161658 77324 161664 77376
rect 161716 77364 161722 77376
rect 167638 77364 167644 77376
rect 161716 77336 167644 77364
rect 161716 77324 161722 77336
rect 167638 77324 167644 77336
rect 167696 77324 167702 77376
rect 169938 77324 169944 77376
rect 169996 77364 170002 77376
rect 170674 77364 170680 77376
rect 169996 77336 170680 77364
rect 169996 77324 170002 77336
rect 170674 77324 170680 77336
rect 170732 77324 170738 77376
rect 176378 77324 176384 77376
rect 176436 77364 176442 77376
rect 177298 77364 177304 77376
rect 176436 77336 177304 77364
rect 176436 77324 176442 77336
rect 177298 77324 177304 77336
rect 177356 77364 177362 77376
rect 179322 77364 179328 77376
rect 177356 77336 179328 77364
rect 177356 77324 177362 77336
rect 179322 77324 179328 77336
rect 179380 77324 179386 77376
rect 132770 77256 132776 77308
rect 132828 77296 132834 77308
rect 132828 77268 133276 77296
rect 132828 77256 132834 77268
rect 105538 77188 105544 77240
rect 105596 77228 105602 77240
rect 105814 77228 105820 77240
rect 105596 77200 105820 77228
rect 105596 77188 105602 77200
rect 105814 77188 105820 77200
rect 105872 77188 105878 77240
rect 124858 77188 124864 77240
rect 124916 77228 124922 77240
rect 125594 77228 125600 77240
rect 124916 77200 125600 77228
rect 124916 77188 124922 77200
rect 125594 77188 125600 77200
rect 125652 77228 125658 77240
rect 133138 77228 133144 77240
rect 125652 77200 133144 77228
rect 125652 77188 125658 77200
rect 133138 77188 133144 77200
rect 133196 77188 133202 77240
rect 133248 77228 133276 77268
rect 162210 77256 162216 77308
rect 162268 77296 162274 77308
rect 177482 77296 177488 77308
rect 162268 77268 177488 77296
rect 162268 77256 162274 77268
rect 177482 77256 177488 77268
rect 177540 77256 177546 77308
rect 137462 77228 137468 77240
rect 133248 77200 137468 77228
rect 137462 77188 137468 77200
rect 137520 77188 137526 77240
rect 159450 77188 159456 77240
rect 159508 77228 159514 77240
rect 161658 77228 161664 77240
rect 159508 77200 161664 77228
rect 159508 77188 159514 77200
rect 161658 77188 161664 77200
rect 161716 77188 161722 77240
rect 172790 77188 172796 77240
rect 172848 77228 172854 77240
rect 205818 77228 205824 77240
rect 172848 77200 205824 77228
rect 172848 77188 172854 77200
rect 205818 77188 205824 77200
rect 205876 77228 205882 77240
rect 206094 77228 206100 77240
rect 205876 77200 206100 77228
rect 205876 77188 205882 77200
rect 206094 77188 206100 77200
rect 206152 77188 206158 77240
rect 122374 77120 122380 77172
rect 122432 77160 122438 77172
rect 144454 77160 144460 77172
rect 122432 77132 144460 77160
rect 122432 77120 122438 77132
rect 144454 77120 144460 77132
rect 144512 77160 144518 77172
rect 145650 77160 145656 77172
rect 144512 77132 145656 77160
rect 144512 77120 144518 77132
rect 145650 77120 145656 77132
rect 145708 77120 145714 77172
rect 156690 77120 156696 77172
rect 156748 77160 156754 77172
rect 156874 77160 156880 77172
rect 156748 77132 156880 77160
rect 156748 77120 156754 77132
rect 156874 77120 156880 77132
rect 156932 77120 156938 77172
rect 161014 77120 161020 77172
rect 161072 77160 161078 77172
rect 191190 77160 191196 77172
rect 161072 77132 191196 77160
rect 161072 77120 161078 77132
rect 191190 77120 191196 77132
rect 191248 77160 191254 77172
rect 191742 77160 191748 77172
rect 191248 77132 191748 77160
rect 191248 77120 191254 77132
rect 191742 77120 191748 77132
rect 191800 77120 191806 77172
rect 118970 77052 118976 77104
rect 119028 77092 119034 77104
rect 119028 77064 142844 77092
rect 119028 77052 119034 77064
rect 108482 76984 108488 77036
rect 108540 77024 108546 77036
rect 108540 76996 133092 77024
rect 108540 76984 108546 76996
rect 105998 76916 106004 76968
rect 106056 76956 106062 76968
rect 130286 76956 130292 76968
rect 106056 76928 130292 76956
rect 106056 76916 106062 76928
rect 130286 76916 130292 76928
rect 130344 76916 130350 76968
rect 132678 76956 132684 76968
rect 130488 76928 132684 76956
rect 118510 76848 118516 76900
rect 118568 76888 118574 76900
rect 130378 76888 130384 76900
rect 118568 76860 130384 76888
rect 118568 76848 118574 76860
rect 130378 76848 130384 76860
rect 130436 76848 130442 76900
rect 106918 76820 106924 76832
rect 103486 76792 106924 76820
rect 72418 76712 72424 76764
rect 72476 76752 72482 76764
rect 103486 76752 103514 76792
rect 106918 76780 106924 76792
rect 106976 76820 106982 76832
rect 130488 76820 130516 76928
rect 132678 76916 132684 76928
rect 132736 76916 132742 76968
rect 133064 76956 133092 76996
rect 133138 76984 133144 77036
rect 133196 77024 133202 77036
rect 141878 77024 141884 77036
rect 133196 76996 141884 77024
rect 133196 76984 133202 76996
rect 141878 76984 141884 76996
rect 141936 76984 141942 77036
rect 142816 77024 142844 77064
rect 147766 77052 147772 77104
rect 147824 77092 147830 77104
rect 147950 77092 147956 77104
rect 147824 77064 147956 77092
rect 147824 77052 147830 77064
rect 147950 77052 147956 77064
rect 148008 77052 148014 77104
rect 159818 77052 159824 77104
rect 159876 77092 159882 77104
rect 189626 77092 189632 77104
rect 159876 77064 189632 77092
rect 159876 77052 159882 77064
rect 189626 77052 189632 77064
rect 189684 77052 189690 77104
rect 152642 77024 152648 77036
rect 142816 76996 152648 77024
rect 152642 76984 152648 76996
rect 152700 77024 152706 77036
rect 152700 76996 153194 77024
rect 152700 76984 152706 76996
rect 133322 76956 133328 76968
rect 133064 76928 133328 76956
rect 133322 76916 133328 76928
rect 133380 76916 133386 76968
rect 144178 76916 144184 76968
rect 144236 76956 144242 76968
rect 151814 76956 151820 76968
rect 144236 76928 151820 76956
rect 144236 76916 144242 76928
rect 151814 76916 151820 76928
rect 151872 76916 151878 76968
rect 133598 76848 133604 76900
rect 133656 76888 133662 76900
rect 133656 76860 138014 76888
rect 133656 76848 133662 76860
rect 106976 76792 130516 76820
rect 106976 76780 106982 76792
rect 134058 76780 134064 76832
rect 134116 76820 134122 76832
rect 136910 76820 136916 76832
rect 134116 76792 136916 76820
rect 134116 76780 134122 76792
rect 136910 76780 136916 76792
rect 136968 76780 136974 76832
rect 137986 76820 138014 76860
rect 149422 76848 149428 76900
rect 149480 76888 149486 76900
rect 149974 76888 149980 76900
rect 149480 76860 149980 76888
rect 149480 76848 149486 76860
rect 149974 76848 149980 76860
rect 150032 76848 150038 76900
rect 148778 76820 148784 76832
rect 137986 76792 148784 76820
rect 148778 76780 148784 76792
rect 148836 76780 148842 76832
rect 72476 76724 103514 76752
rect 72476 76712 72482 76724
rect 119430 76712 119436 76764
rect 119488 76752 119494 76764
rect 148594 76752 148600 76764
rect 119488 76724 148600 76752
rect 119488 76712 119494 76724
rect 148594 76712 148600 76724
rect 148652 76712 148658 76764
rect 153166 76752 153194 76996
rect 177942 76984 177948 77036
rect 178000 77024 178006 77036
rect 205910 77024 205916 77036
rect 178000 76996 205916 77024
rect 178000 76984 178006 76996
rect 205910 76984 205916 76996
rect 205968 76984 205974 77036
rect 155494 76916 155500 76968
rect 155552 76956 155558 76968
rect 179322 76956 179328 76968
rect 155552 76928 179328 76956
rect 155552 76916 155558 76928
rect 179322 76916 179328 76928
rect 179380 76916 179386 76968
rect 170214 76848 170220 76900
rect 170272 76888 170278 76900
rect 170582 76888 170588 76900
rect 170272 76860 170588 76888
rect 170272 76848 170278 76860
rect 170582 76848 170588 76860
rect 170640 76888 170646 76900
rect 192570 76888 192576 76900
rect 170640 76860 192576 76888
rect 170640 76848 170646 76860
rect 192570 76848 192576 76860
rect 192628 76848 192634 76900
rect 170674 76780 170680 76832
rect 170732 76820 170738 76832
rect 192754 76820 192760 76832
rect 170732 76792 192760 76820
rect 170732 76780 170738 76792
rect 192754 76780 192760 76792
rect 192812 76780 192818 76832
rect 260834 76752 260840 76764
rect 153166 76724 260840 76752
rect 260834 76712 260840 76724
rect 260892 76712 260898 76764
rect 64138 76644 64144 76696
rect 64196 76684 64202 76696
rect 105998 76684 106004 76696
rect 64196 76656 106004 76684
rect 64196 76644 64202 76656
rect 105998 76644 106004 76656
rect 106056 76644 106062 76696
rect 117406 76644 117412 76696
rect 117464 76684 117470 76696
rect 132770 76684 132776 76696
rect 117464 76656 132776 76684
rect 117464 76644 117470 76656
rect 132770 76644 132776 76656
rect 132828 76644 132834 76696
rect 134518 76644 134524 76696
rect 134576 76684 134582 76696
rect 139026 76684 139032 76696
rect 134576 76656 139032 76684
rect 134576 76644 134582 76656
rect 139026 76644 139032 76656
rect 139084 76644 139090 76696
rect 143534 76644 143540 76696
rect 143592 76684 143598 76696
rect 144086 76684 144092 76696
rect 143592 76656 144092 76684
rect 143592 76644 143598 76656
rect 144086 76644 144092 76656
rect 144144 76644 144150 76696
rect 148318 76644 148324 76696
rect 148376 76684 148382 76696
rect 148686 76684 148692 76696
rect 148376 76656 148692 76684
rect 148376 76644 148382 76656
rect 148686 76644 148692 76656
rect 148744 76644 148750 76696
rect 149330 76644 149336 76696
rect 149388 76684 149394 76696
rect 149388 76656 161474 76684
rect 149388 76644 149394 76656
rect 52454 76576 52460 76628
rect 52512 76616 52518 76628
rect 135806 76616 135812 76628
rect 52512 76588 135812 76616
rect 52512 76576 52518 76588
rect 135806 76576 135812 76588
rect 135864 76576 135870 76628
rect 149606 76576 149612 76628
rect 149664 76616 149670 76628
rect 150250 76616 150256 76628
rect 149664 76588 150256 76616
rect 149664 76576 149670 76588
rect 150250 76576 150256 76588
rect 150308 76576 150314 76628
rect 161446 76616 161474 76656
rect 161750 76644 161756 76696
rect 161808 76684 161814 76696
rect 161934 76684 161940 76696
rect 161808 76656 161940 76684
rect 161808 76644 161814 76656
rect 161934 76644 161940 76656
rect 161992 76644 161998 76696
rect 162854 76644 162860 76696
rect 162912 76684 162918 76696
rect 163038 76684 163044 76696
rect 162912 76656 163044 76684
rect 162912 76644 162918 76656
rect 163038 76644 163044 76656
rect 163096 76644 163102 76696
rect 167178 76644 167184 76696
rect 167236 76684 167242 76696
rect 169110 76684 169116 76696
rect 167236 76656 169116 76684
rect 167236 76644 167242 76656
rect 169110 76644 169116 76656
rect 169168 76644 169174 76696
rect 170858 76644 170864 76696
rect 170916 76684 170922 76696
rect 189534 76684 189540 76696
rect 170916 76656 189540 76684
rect 170916 76644 170922 76656
rect 189534 76644 189540 76656
rect 189592 76644 189598 76696
rect 189626 76644 189632 76696
rect 189684 76684 189690 76696
rect 353294 76684 353300 76696
rect 189684 76656 353300 76684
rect 189684 76644 189690 76656
rect 353294 76644 353300 76656
rect 353352 76644 353358 76696
rect 181438 76616 181444 76628
rect 161446 76588 181444 76616
rect 181438 76576 181444 76588
rect 181496 76576 181502 76628
rect 191742 76576 191748 76628
rect 191800 76616 191806 76628
rect 367094 76616 367100 76628
rect 191800 76588 367100 76616
rect 191800 76576 191806 76588
rect 367094 76576 367100 76588
rect 367152 76576 367158 76628
rect 35894 76508 35900 76560
rect 35952 76548 35958 76560
rect 135254 76548 135260 76560
rect 35952 76520 135260 76548
rect 35952 76508 35958 76520
rect 135254 76508 135260 76520
rect 135312 76508 135318 76560
rect 151262 76508 151268 76560
rect 151320 76548 151326 76560
rect 203702 76548 203708 76560
rect 151320 76520 203708 76548
rect 151320 76508 151326 76520
rect 203702 76508 203708 76520
rect 203760 76508 203766 76560
rect 205818 76508 205824 76560
rect 205876 76548 205882 76560
rect 509878 76548 509884 76560
rect 205876 76520 509884 76548
rect 205876 76508 205882 76520
rect 509878 76508 509884 76520
rect 509936 76508 509942 76560
rect 126238 76440 126244 76492
rect 126296 76480 126302 76492
rect 133138 76480 133144 76492
rect 126296 76452 133144 76480
rect 126296 76440 126302 76452
rect 133138 76440 133144 76452
rect 133196 76440 133202 76492
rect 133322 76440 133328 76492
rect 133380 76480 133386 76492
rect 140406 76480 140412 76492
rect 133380 76452 140412 76480
rect 133380 76440 133386 76452
rect 140406 76440 140412 76452
rect 140464 76440 140470 76492
rect 161750 76440 161756 76492
rect 161808 76480 161814 76492
rect 162394 76480 162400 76492
rect 161808 76452 162400 76480
rect 161808 76440 161814 76452
rect 162394 76440 162400 76452
rect 162452 76440 162458 76492
rect 162854 76440 162860 76492
rect 162912 76480 162918 76492
rect 164234 76480 164240 76492
rect 162912 76452 164240 76480
rect 162912 76440 162918 76452
rect 164234 76440 164240 76452
rect 164292 76440 164298 76492
rect 168558 76440 168564 76492
rect 168616 76480 168622 76492
rect 168742 76480 168748 76492
rect 168616 76452 168748 76480
rect 168616 76440 168622 76452
rect 168742 76440 168748 76452
rect 168800 76440 168806 76492
rect 169018 76440 169024 76492
rect 169076 76480 169082 76492
rect 178678 76480 178684 76492
rect 169076 76452 178684 76480
rect 169076 76440 169082 76452
rect 178678 76440 178684 76452
rect 178736 76440 178742 76492
rect 112438 76372 112444 76424
rect 112496 76412 112502 76424
rect 146662 76412 146668 76424
rect 112496 76384 146668 76412
rect 112496 76372 112502 76384
rect 146662 76372 146668 76384
rect 146720 76412 146726 76424
rect 153930 76412 153936 76424
rect 146720 76384 153936 76412
rect 146720 76372 146726 76384
rect 153930 76372 153936 76384
rect 153988 76372 153994 76424
rect 160830 76372 160836 76424
rect 160888 76412 160894 76424
rect 161290 76412 161296 76424
rect 160888 76384 161296 76412
rect 160888 76372 160894 76384
rect 161290 76372 161296 76384
rect 161348 76372 161354 76424
rect 168834 76372 168840 76424
rect 168892 76412 168898 76424
rect 169202 76412 169208 76424
rect 168892 76384 169208 76412
rect 168892 76372 168898 76384
rect 169202 76372 169208 76384
rect 169260 76372 169266 76424
rect 105538 76304 105544 76356
rect 105596 76344 105602 76356
rect 105596 76316 122834 76344
rect 105596 76304 105602 76316
rect 122806 76276 122834 76316
rect 132770 76304 132776 76356
rect 132828 76344 132834 76356
rect 141050 76344 141056 76356
rect 132828 76316 141056 76344
rect 132828 76304 132834 76316
rect 141050 76304 141056 76316
rect 141108 76304 141114 76356
rect 171962 76304 171968 76356
rect 172020 76344 172026 76356
rect 189718 76344 189724 76356
rect 172020 76316 189724 76344
rect 172020 76304 172026 76316
rect 189718 76304 189724 76316
rect 189776 76304 189782 76356
rect 140130 76276 140136 76288
rect 122806 76248 140136 76276
rect 140130 76236 140136 76248
rect 140188 76236 140194 76288
rect 133138 76168 133144 76220
rect 133196 76208 133202 76220
rect 141694 76208 141700 76220
rect 133196 76180 141700 76208
rect 133196 76168 133202 76180
rect 141694 76168 141700 76180
rect 141752 76168 141758 76220
rect 164234 76168 164240 76220
rect 164292 76208 164298 76220
rect 165798 76208 165804 76220
rect 164292 76180 165804 76208
rect 164292 76168 164298 76180
rect 165798 76168 165804 76180
rect 165856 76168 165862 76220
rect 164602 76032 164608 76084
rect 164660 76072 164666 76084
rect 164878 76072 164884 76084
rect 164660 76044 164884 76072
rect 164660 76032 164666 76044
rect 164878 76032 164884 76044
rect 164936 76032 164942 76084
rect 172698 76032 172704 76084
rect 172756 76072 172762 76084
rect 173618 76072 173624 76084
rect 172756 76044 173624 76072
rect 172756 76032 172762 76044
rect 173618 76032 173624 76044
rect 173676 76032 173682 76084
rect 158622 75964 158628 76016
rect 158680 76004 158686 76016
rect 180058 76004 180064 76016
rect 158680 75976 180064 76004
rect 158680 75964 158686 75976
rect 180058 75964 180064 75976
rect 180116 76004 180122 76016
rect 289814 76004 289820 76016
rect 180116 75976 289820 76004
rect 180116 75964 180122 75976
rect 289814 75964 289820 75976
rect 289872 75964 289878 76016
rect 110708 75908 111196 75936
rect 104894 75828 104900 75880
rect 104952 75868 104958 75880
rect 110708 75868 110736 75908
rect 104952 75840 110736 75868
rect 104952 75828 104958 75840
rect 110782 75828 110788 75880
rect 110840 75868 110846 75880
rect 111058 75868 111064 75880
rect 110840 75840 111064 75868
rect 110840 75828 110846 75840
rect 111058 75828 111064 75840
rect 111116 75828 111122 75880
rect 111168 75868 111196 75908
rect 146018 75896 146024 75948
rect 146076 75936 146082 75948
rect 146938 75936 146944 75948
rect 146076 75908 146944 75936
rect 146076 75896 146082 75908
rect 146938 75896 146944 75908
rect 146996 75896 147002 75948
rect 164510 75896 164516 75948
rect 164568 75936 164574 75948
rect 165154 75936 165160 75948
rect 164568 75908 165160 75936
rect 164568 75896 164574 75908
rect 165154 75896 165160 75908
rect 165212 75896 165218 75948
rect 167086 75896 167092 75948
rect 167144 75936 167150 75948
rect 167730 75936 167736 75948
rect 167144 75908 167736 75936
rect 167144 75896 167150 75908
rect 167730 75896 167736 75908
rect 167788 75896 167794 75948
rect 171962 75896 171968 75948
rect 172020 75936 172026 75948
rect 172146 75936 172152 75948
rect 172020 75908 172152 75936
rect 172020 75896 172026 75908
rect 172146 75896 172152 75908
rect 172204 75896 172210 75948
rect 179322 75896 179328 75948
rect 179380 75936 179386 75948
rect 296714 75936 296720 75948
rect 179380 75908 296720 75936
rect 179380 75896 179386 75908
rect 296714 75896 296720 75908
rect 296772 75896 296778 75948
rect 139394 75868 139400 75880
rect 111168 75840 139400 75868
rect 139394 75828 139400 75840
rect 139452 75828 139458 75880
rect 144454 75828 144460 75880
rect 144512 75868 144518 75880
rect 151078 75868 151084 75880
rect 144512 75840 151084 75868
rect 144512 75828 144518 75840
rect 151078 75828 151084 75840
rect 151136 75828 151142 75880
rect 163590 75828 163596 75880
rect 163648 75868 163654 75880
rect 163866 75868 163872 75880
rect 163648 75840 163872 75868
rect 163648 75828 163654 75840
rect 163866 75828 163872 75840
rect 163924 75868 163930 75880
rect 198458 75868 198464 75880
rect 163924 75840 198464 75868
rect 163924 75828 163930 75840
rect 198458 75828 198464 75840
rect 198516 75828 198522 75880
rect 107010 75760 107016 75812
rect 107068 75800 107074 75812
rect 138014 75800 138020 75812
rect 107068 75772 138020 75800
rect 107068 75760 107074 75772
rect 138014 75760 138020 75772
rect 138072 75760 138078 75812
rect 164418 75760 164424 75812
rect 164476 75800 164482 75812
rect 165430 75800 165436 75812
rect 164476 75772 165436 75800
rect 164476 75760 164482 75772
rect 165430 75760 165436 75772
rect 165488 75760 165494 75812
rect 165798 75760 165804 75812
rect 165856 75800 165862 75812
rect 166074 75800 166080 75812
rect 165856 75772 166080 75800
rect 165856 75760 165862 75772
rect 166074 75760 166080 75772
rect 166132 75760 166138 75812
rect 166902 75760 166908 75812
rect 166960 75800 166966 75812
rect 167178 75800 167184 75812
rect 166960 75772 167184 75800
rect 166960 75760 166966 75772
rect 167178 75760 167184 75772
rect 167236 75760 167242 75812
rect 171410 75760 171416 75812
rect 171468 75800 171474 75812
rect 171962 75800 171968 75812
rect 171468 75772 171968 75800
rect 171468 75760 171474 75772
rect 171962 75760 171968 75772
rect 172020 75760 172026 75812
rect 187970 75800 187976 75812
rect 172670 75772 187976 75800
rect 115382 75692 115388 75744
rect 115440 75732 115446 75744
rect 146386 75732 146392 75744
rect 115440 75704 146392 75732
rect 115440 75692 115446 75704
rect 146386 75692 146392 75704
rect 146444 75732 146450 75744
rect 154298 75732 154304 75744
rect 146444 75704 154304 75732
rect 146444 75692 146450 75704
rect 154298 75692 154304 75704
rect 154356 75692 154362 75744
rect 163130 75692 163136 75744
rect 163188 75732 163194 75744
rect 166258 75732 166264 75744
rect 163188 75704 166264 75732
rect 163188 75692 163194 75704
rect 166258 75692 166264 75704
rect 166316 75692 166322 75744
rect 170398 75692 170404 75744
rect 170456 75732 170462 75744
rect 171042 75732 171048 75744
rect 170456 75704 171048 75732
rect 170456 75692 170462 75704
rect 171042 75692 171048 75704
rect 171100 75732 171106 75744
rect 172670 75732 172698 75772
rect 187970 75760 187976 75772
rect 188028 75760 188034 75812
rect 171100 75704 172698 75732
rect 171100 75692 171106 75704
rect 178494 75692 178500 75744
rect 178552 75732 178558 75744
rect 183554 75732 183560 75744
rect 178552 75704 183560 75732
rect 178552 75692 178558 75704
rect 183554 75692 183560 75704
rect 183612 75692 183618 75744
rect 111058 75624 111064 75676
rect 111116 75664 111122 75676
rect 139946 75664 139952 75676
rect 111116 75636 139952 75664
rect 111116 75624 111122 75636
rect 139946 75624 139952 75636
rect 140004 75624 140010 75676
rect 146754 75624 146760 75676
rect 146812 75664 146818 75676
rect 182818 75664 182824 75676
rect 146812 75636 182824 75664
rect 146812 75624 146818 75636
rect 182818 75624 182824 75636
rect 182876 75624 182882 75676
rect 108666 75556 108672 75608
rect 108724 75596 108730 75608
rect 135438 75596 135444 75608
rect 108724 75568 135444 75596
rect 108724 75556 108730 75568
rect 135438 75556 135444 75568
rect 135496 75556 135502 75608
rect 153930 75556 153936 75608
rect 153988 75596 153994 75608
rect 187694 75596 187700 75608
rect 153988 75568 187700 75596
rect 153988 75556 153994 75568
rect 187694 75556 187700 75568
rect 187752 75556 187758 75608
rect 115198 75488 115204 75540
rect 115256 75528 115262 75540
rect 117406 75528 117412 75540
rect 115256 75500 117412 75528
rect 115256 75488 115262 75500
rect 117406 75488 117412 75500
rect 117464 75488 117470 75540
rect 121270 75488 121276 75540
rect 121328 75528 121334 75540
rect 146570 75528 146576 75540
rect 121328 75500 146576 75528
rect 121328 75488 121334 75500
rect 146570 75488 146576 75500
rect 146628 75528 146634 75540
rect 147950 75528 147956 75540
rect 146628 75500 147956 75528
rect 146628 75488 146634 75500
rect 147950 75488 147956 75500
rect 148008 75488 148014 75540
rect 148042 75488 148048 75540
rect 148100 75528 148106 75540
rect 201494 75528 201500 75540
rect 148100 75500 201500 75528
rect 148100 75488 148106 75500
rect 201494 75488 201500 75500
rect 201552 75488 201558 75540
rect 122558 75420 122564 75472
rect 122616 75460 122622 75472
rect 145190 75460 145196 75472
rect 122616 75432 145196 75460
rect 122616 75420 122622 75432
rect 145190 75420 145196 75432
rect 145248 75420 145254 75472
rect 150342 75420 150348 75472
rect 150400 75460 150406 75472
rect 216674 75460 216680 75472
rect 150400 75432 216680 75460
rect 150400 75420 150406 75432
rect 216674 75420 216680 75432
rect 216732 75420 216738 75472
rect 81434 75352 81440 75404
rect 81492 75392 81498 75404
rect 138658 75392 138664 75404
rect 81492 75364 138664 75392
rect 81492 75352 81498 75364
rect 138658 75352 138664 75364
rect 138716 75352 138722 75404
rect 166350 75352 166356 75404
rect 166408 75392 166414 75404
rect 166902 75392 166908 75404
rect 166408 75364 166908 75392
rect 166408 75352 166414 75364
rect 166902 75352 166908 75364
rect 166960 75352 166966 75404
rect 172974 75352 172980 75404
rect 173032 75392 173038 75404
rect 480898 75392 480904 75404
rect 173032 75364 480904 75392
rect 173032 75352 173038 75364
rect 480898 75352 480904 75364
rect 480956 75352 480962 75404
rect 67634 75284 67640 75336
rect 67692 75324 67698 75336
rect 137646 75324 137652 75336
rect 67692 75296 137652 75324
rect 67692 75284 67698 75296
rect 137646 75284 137652 75296
rect 137704 75284 137710 75336
rect 145098 75284 145104 75336
rect 145156 75324 145162 75336
rect 145742 75324 145748 75336
rect 145156 75296 145748 75324
rect 145156 75284 145162 75296
rect 145742 75284 145748 75296
rect 145800 75284 145806 75336
rect 172238 75284 172244 75336
rect 172296 75324 172302 75336
rect 506474 75324 506480 75336
rect 172296 75296 506480 75324
rect 172296 75284 172302 75296
rect 506474 75284 506480 75296
rect 506532 75284 506538 75336
rect 22738 75216 22744 75268
rect 22796 75256 22802 75268
rect 132402 75256 132408 75268
rect 22796 75228 132408 75256
rect 22796 75216 22802 75228
rect 132402 75216 132408 75228
rect 132460 75216 132466 75268
rect 135806 75216 135812 75268
rect 135864 75256 135870 75268
rect 136358 75256 136364 75268
rect 135864 75228 136364 75256
rect 135864 75216 135870 75228
rect 136358 75216 136364 75228
rect 136416 75216 136422 75268
rect 139486 75216 139492 75268
rect 139544 75256 139550 75268
rect 140314 75256 140320 75268
rect 139544 75228 140320 75256
rect 139544 75216 139550 75228
rect 140314 75216 140320 75228
rect 140372 75216 140378 75268
rect 153194 75216 153200 75268
rect 153252 75256 153258 75268
rect 153838 75256 153844 75268
rect 153252 75228 153844 75256
rect 153252 75216 153258 75228
rect 153838 75216 153844 75228
rect 153896 75216 153902 75268
rect 158898 75216 158904 75268
rect 158956 75256 158962 75268
rect 159174 75256 159180 75268
rect 158956 75228 159180 75256
rect 158956 75216 158962 75228
rect 159174 75216 159180 75228
rect 159232 75216 159238 75268
rect 172330 75216 172336 75268
rect 172388 75256 172394 75268
rect 511258 75256 511264 75268
rect 172388 75228 511264 75256
rect 172388 75216 172394 75228
rect 511258 75216 511264 75228
rect 511316 75216 511322 75268
rect 7558 75148 7564 75200
rect 7616 75188 7622 75200
rect 120074 75188 120080 75200
rect 7616 75160 120080 75188
rect 7616 75148 7622 75160
rect 120074 75148 120080 75160
rect 120132 75148 120138 75200
rect 122282 75148 122288 75200
rect 122340 75188 122346 75200
rect 145558 75188 145564 75200
rect 122340 75160 145564 75188
rect 122340 75148 122346 75160
rect 145558 75148 145564 75160
rect 145616 75148 145622 75200
rect 168006 75148 168012 75200
rect 168064 75188 168070 75200
rect 168064 75160 171134 75188
rect 168064 75148 168070 75160
rect 130010 75080 130016 75132
rect 130068 75120 130074 75132
rect 131022 75120 131028 75132
rect 130068 75092 131028 75120
rect 130068 75080 130074 75092
rect 131022 75080 131028 75092
rect 131080 75080 131086 75132
rect 162670 75080 162676 75132
rect 162728 75120 162734 75132
rect 164786 75120 164792 75132
rect 162728 75092 164792 75120
rect 162728 75080 162734 75092
rect 164786 75080 164792 75092
rect 164844 75080 164850 75132
rect 168742 75080 168748 75132
rect 168800 75120 168806 75132
rect 169294 75120 169300 75132
rect 168800 75092 169300 75120
rect 168800 75080 168806 75092
rect 169294 75080 169300 75092
rect 169352 75080 169358 75132
rect 171106 75120 171134 75160
rect 178034 75148 178040 75200
rect 178092 75188 178098 75200
rect 549254 75188 549260 75200
rect 178092 75160 549260 75188
rect 178092 75148 178098 75160
rect 549254 75148 549260 75160
rect 549312 75148 549318 75200
rect 171106 75092 176654 75120
rect 154114 75012 154120 75064
rect 154172 75052 154178 75064
rect 154390 75052 154396 75064
rect 154172 75024 154396 75052
rect 154172 75012 154178 75024
rect 154390 75012 154396 75024
rect 154448 75012 154454 75064
rect 176626 75052 176654 75092
rect 176838 75080 176844 75132
rect 176896 75120 176902 75132
rect 177114 75120 177120 75132
rect 176896 75092 177120 75120
rect 176896 75080 176902 75092
rect 177114 75080 177120 75092
rect 177172 75080 177178 75132
rect 177758 75080 177764 75132
rect 177816 75120 177822 75132
rect 177816 75092 186314 75120
rect 177816 75080 177822 75092
rect 180058 75052 180064 75064
rect 176626 75024 180064 75052
rect 180058 75012 180064 75024
rect 180116 75012 180122 75064
rect 186286 75052 186314 75092
rect 205726 75052 205732 75064
rect 186286 75024 205732 75052
rect 205726 75012 205732 75024
rect 205784 75012 205790 75064
rect 154298 74944 154304 74996
rect 154356 74984 154362 74996
rect 180794 74984 180800 74996
rect 154356 74956 180800 74984
rect 154356 74944 154362 74956
rect 180794 74944 180800 74956
rect 180852 74944 180858 74996
rect 135438 74876 135444 74928
rect 135496 74916 135502 74928
rect 136542 74916 136548 74928
rect 135496 74888 136548 74916
rect 135496 74876 135502 74888
rect 136542 74876 136548 74888
rect 136600 74876 136606 74928
rect 177022 74876 177028 74928
rect 177080 74916 177086 74928
rect 177482 74916 177488 74928
rect 177080 74888 177488 74916
rect 177080 74876 177086 74888
rect 177482 74876 177488 74888
rect 177540 74876 177546 74928
rect 132954 74740 132960 74792
rect 133012 74780 133018 74792
rect 133506 74780 133512 74792
rect 133012 74752 133512 74780
rect 133012 74740 133018 74752
rect 133506 74740 133512 74752
rect 133564 74740 133570 74792
rect 143994 74576 144000 74588
rect 139366 74548 144000 74576
rect 109954 74468 109960 74520
rect 110012 74508 110018 74520
rect 139366 74508 139394 74548
rect 143994 74536 144000 74548
rect 144052 74536 144058 74588
rect 175826 74536 175832 74588
rect 175884 74576 175890 74588
rect 176102 74576 176108 74588
rect 175884 74548 176108 74576
rect 175884 74536 175890 74548
rect 176102 74536 176108 74548
rect 176160 74536 176166 74588
rect 110012 74480 139394 74508
rect 110012 74468 110018 74480
rect 142246 74468 142252 74520
rect 142304 74508 142310 74520
rect 143166 74508 143172 74520
rect 142304 74480 143172 74508
rect 142304 74468 142310 74480
rect 143166 74468 143172 74480
rect 143224 74468 143230 74520
rect 153286 74468 153292 74520
rect 153344 74508 153350 74520
rect 154022 74508 154028 74520
rect 153344 74480 154028 74508
rect 153344 74468 153350 74480
rect 154022 74468 154028 74480
rect 154080 74468 154086 74520
rect 166902 74468 166908 74520
rect 166960 74508 166966 74520
rect 200942 74508 200948 74520
rect 166960 74480 200948 74508
rect 166960 74468 166966 74480
rect 200942 74468 200948 74480
rect 201000 74468 201006 74520
rect 110046 74400 110052 74452
rect 110104 74440 110110 74452
rect 144638 74440 144644 74452
rect 110104 74412 144644 74440
rect 110104 74400 110110 74412
rect 144638 74400 144644 74412
rect 144696 74400 144702 74452
rect 153378 74400 153384 74452
rect 153436 74440 153442 74452
rect 188614 74440 188620 74452
rect 153436 74412 188620 74440
rect 153436 74400 153442 74412
rect 188614 74400 188620 74412
rect 188672 74440 188678 74452
rect 269114 74440 269120 74452
rect 188672 74412 269120 74440
rect 188672 74400 188678 74412
rect 269114 74400 269120 74412
rect 269172 74400 269178 74452
rect 112898 74332 112904 74384
rect 112956 74372 112962 74384
rect 112956 74344 143120 74372
rect 112956 74332 112962 74344
rect 111518 74264 111524 74316
rect 111576 74304 111582 74316
rect 141510 74304 141516 74316
rect 111576 74276 141516 74304
rect 111576 74264 111582 74276
rect 141510 74264 141516 74276
rect 141568 74264 141574 74316
rect 143092 74304 143120 74344
rect 143166 74332 143172 74384
rect 143224 74372 143230 74384
rect 143442 74372 143448 74384
rect 143224 74344 143448 74372
rect 143224 74332 143230 74344
rect 143442 74332 143448 74344
rect 143500 74332 143506 74384
rect 171502 74332 171508 74384
rect 171560 74372 171566 74384
rect 172146 74372 172152 74384
rect 171560 74344 172152 74372
rect 171560 74332 171566 74344
rect 172146 74332 172152 74344
rect 172204 74332 172210 74384
rect 172882 74332 172888 74384
rect 172940 74372 172946 74384
rect 173526 74372 173532 74384
rect 172940 74344 173532 74372
rect 172940 74332 172946 74344
rect 173526 74332 173532 74344
rect 173584 74372 173590 74384
rect 198274 74372 198280 74384
rect 173584 74344 198280 74372
rect 173584 74332 173590 74344
rect 198274 74332 198280 74344
rect 198332 74332 198338 74384
rect 144914 74304 144920 74316
rect 143092 74276 144920 74304
rect 144914 74264 144920 74276
rect 144972 74264 144978 74316
rect 172514 74264 172520 74316
rect 172572 74304 172578 74316
rect 173434 74304 173440 74316
rect 172572 74276 173440 74304
rect 172572 74264 172578 74276
rect 173434 74264 173440 74276
rect 173492 74304 173498 74316
rect 196986 74304 196992 74316
rect 173492 74276 196992 74304
rect 173492 74264 173498 74276
rect 196986 74264 196992 74276
rect 197044 74264 197050 74316
rect 111426 74196 111432 74248
rect 111484 74236 111490 74248
rect 143902 74236 143908 74248
rect 111484 74208 143908 74236
rect 111484 74196 111490 74208
rect 143902 74196 143908 74208
rect 143960 74236 143966 74248
rect 147122 74236 147128 74248
rect 143960 74208 147128 74236
rect 143960 74196 143966 74208
rect 147122 74196 147128 74208
rect 147180 74196 147186 74248
rect 150986 74196 150992 74248
rect 151044 74236 151050 74248
rect 237374 74236 237380 74248
rect 151044 74208 237380 74236
rect 151044 74196 151050 74208
rect 237374 74196 237380 74208
rect 237432 74196 237438 74248
rect 100202 74128 100208 74180
rect 100260 74168 100266 74180
rect 133782 74168 133788 74180
rect 100260 74140 133788 74168
rect 100260 74128 100266 74140
rect 133782 74128 133788 74140
rect 133840 74128 133846 74180
rect 141510 74128 141516 74180
rect 141568 74168 141574 74180
rect 144546 74168 144552 74180
rect 141568 74140 144552 74168
rect 141568 74128 141574 74140
rect 144546 74128 144552 74140
rect 144604 74128 144610 74180
rect 152366 74128 152372 74180
rect 152424 74168 152430 74180
rect 255314 74168 255320 74180
rect 152424 74140 255320 74168
rect 152424 74128 152430 74140
rect 255314 74128 255320 74140
rect 255372 74128 255378 74180
rect 104158 74060 104164 74112
rect 104216 74100 104222 74112
rect 135530 74100 135536 74112
rect 104216 74072 135536 74100
rect 104216 74060 104222 74072
rect 135530 74060 135536 74072
rect 135588 74060 135594 74112
rect 153470 74060 153476 74112
rect 153528 74100 153534 74112
rect 284294 74100 284300 74112
rect 153528 74072 284300 74100
rect 153528 74060 153534 74072
rect 284294 74060 284300 74072
rect 284352 74060 284358 74112
rect 93854 73992 93860 74044
rect 93912 74032 93918 74044
rect 104894 74032 104900 74044
rect 93912 74004 104900 74032
rect 93912 73992 93918 74004
rect 104894 73992 104900 74004
rect 104952 73992 104958 74044
rect 123202 73992 123208 74044
rect 123260 74032 123266 74044
rect 153286 74032 153292 74044
rect 123260 74004 153292 74032
rect 123260 73992 123266 74004
rect 153286 73992 153292 74004
rect 153344 73992 153350 74044
rect 155586 73992 155592 74044
rect 155644 74032 155650 74044
rect 297358 74032 297364 74044
rect 155644 74004 297364 74032
rect 155644 73992 155650 74004
rect 297358 73992 297364 74004
rect 297416 73992 297422 74044
rect 104250 73924 104256 73976
rect 104308 73964 104314 73976
rect 134150 73964 134156 73976
rect 104308 73936 134156 73964
rect 104308 73924 104314 73936
rect 134150 73924 134156 73936
rect 134208 73964 134214 73976
rect 134610 73964 134616 73976
rect 134208 73936 134616 73964
rect 134208 73924 134214 73936
rect 134610 73924 134616 73936
rect 134668 73924 134674 73976
rect 161658 73924 161664 73976
rect 161716 73964 161722 73976
rect 347774 73964 347780 73976
rect 161716 73936 347780 73964
rect 161716 73924 161722 73936
rect 347774 73924 347780 73936
rect 347832 73924 347838 73976
rect 54478 73856 54484 73908
rect 54536 73896 54542 73908
rect 107562 73896 107568 73908
rect 54536 73868 107568 73896
rect 54536 73856 54542 73868
rect 107562 73856 107568 73868
rect 107620 73856 107626 73908
rect 112806 73856 112812 73908
rect 112864 73896 112870 73908
rect 142246 73896 142252 73908
rect 112864 73868 142252 73896
rect 112864 73856 112870 73868
rect 142246 73856 142252 73868
rect 142304 73856 142310 73908
rect 152734 73856 152740 73908
rect 152792 73896 152798 73908
rect 261478 73896 261484 73908
rect 152792 73868 261484 73896
rect 152792 73856 152798 73868
rect 261478 73856 261484 73868
rect 261536 73856 261542 73908
rect 269758 73856 269764 73908
rect 269816 73896 269822 73908
rect 465166 73896 465172 73908
rect 269816 73868 465172 73896
rect 269816 73856 269822 73868
rect 465166 73856 465172 73868
rect 465224 73856 465230 73908
rect 21358 73788 21364 73840
rect 21416 73828 21422 73840
rect 100202 73828 100208 73840
rect 21416 73800 100208 73828
rect 21416 73788 21422 73800
rect 100202 73788 100208 73800
rect 100260 73788 100266 73840
rect 112990 73788 112996 73840
rect 113048 73828 113054 73840
rect 142522 73828 142528 73840
rect 113048 73800 142528 73828
rect 113048 73788 113054 73800
rect 142522 73788 142528 73800
rect 142580 73788 142586 73840
rect 151722 73788 151728 73840
rect 151780 73828 151786 73840
rect 248414 73828 248420 73840
rect 151780 73800 248420 73828
rect 151780 73788 151786 73800
rect 248414 73788 248420 73800
rect 248472 73788 248478 73840
rect 253198 73788 253204 73840
rect 253256 73828 253262 73840
rect 449894 73828 449900 73840
rect 253256 73800 449900 73828
rect 253256 73788 253262 73800
rect 449894 73788 449900 73800
rect 449952 73788 449958 73840
rect 114186 73720 114192 73772
rect 114244 73760 114250 73772
rect 142982 73760 142988 73772
rect 114244 73732 142988 73760
rect 114244 73720 114250 73732
rect 142982 73720 142988 73732
rect 143040 73720 143046 73772
rect 155034 73720 155040 73772
rect 155092 73760 155098 73772
rect 155678 73760 155684 73772
rect 155092 73732 155684 73760
rect 155092 73720 155098 73732
rect 155678 73720 155684 73732
rect 155736 73720 155742 73772
rect 172514 73720 172520 73772
rect 172572 73760 172578 73772
rect 173342 73760 173348 73772
rect 172572 73732 173348 73760
rect 172572 73720 172578 73732
rect 173342 73720 173348 73732
rect 173400 73720 173406 73772
rect 192386 73760 192392 73772
rect 176626 73732 192392 73760
rect 107562 73652 107568 73704
rect 107620 73692 107626 73704
rect 136450 73692 136456 73704
rect 107620 73664 136456 73692
rect 107620 73652 107626 73664
rect 136450 73652 136456 73664
rect 136508 73652 136514 73704
rect 172146 73652 172152 73704
rect 172204 73692 172210 73704
rect 176626 73692 176654 73732
rect 192386 73720 192392 73732
rect 192444 73720 192450 73772
rect 172204 73664 176654 73692
rect 172204 73652 172210 73664
rect 104250 73312 104256 73364
rect 104308 73352 104314 73364
rect 104618 73352 104624 73364
rect 104308 73324 104624 73352
rect 104308 73312 104314 73324
rect 104618 73312 104624 73324
rect 104676 73312 104682 73364
rect 111334 73176 111340 73228
rect 111392 73216 111398 73228
rect 114554 73216 114560 73228
rect 111392 73188 114560 73216
rect 111392 73176 111398 73188
rect 114554 73176 114560 73188
rect 114612 73216 114618 73228
rect 115842 73216 115848 73228
rect 114612 73188 115848 73216
rect 114612 73176 114618 73188
rect 115842 73176 115848 73188
rect 115900 73176 115906 73228
rect 110230 73108 110236 73160
rect 110288 73148 110294 73160
rect 144086 73148 144092 73160
rect 110288 73120 144092 73148
rect 110288 73108 110294 73120
rect 144086 73108 144092 73120
rect 144144 73108 144150 73160
rect 157334 73108 157340 73160
rect 157392 73148 157398 73160
rect 158254 73148 158260 73160
rect 157392 73120 158260 73148
rect 157392 73108 157398 73120
rect 158254 73108 158260 73120
rect 158312 73108 158318 73160
rect 160370 73108 160376 73160
rect 160428 73148 160434 73160
rect 161106 73148 161112 73160
rect 160428 73120 161112 73148
rect 160428 73108 160434 73120
rect 161106 73108 161112 73120
rect 161164 73108 161170 73160
rect 167822 73108 167828 73160
rect 167880 73148 167886 73160
rect 168006 73148 168012 73160
rect 167880 73120 168012 73148
rect 167880 73108 167886 73120
rect 168006 73108 168012 73120
rect 168064 73148 168070 73160
rect 202322 73148 202328 73160
rect 168064 73120 202328 73148
rect 168064 73108 168070 73120
rect 202322 73108 202328 73120
rect 202380 73108 202386 73160
rect 327718 73108 327724 73160
rect 327776 73148 327782 73160
rect 580166 73148 580172 73160
rect 327776 73120 580172 73148
rect 327776 73108 327782 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 123754 73040 123760 73092
rect 123812 73080 123818 73092
rect 149330 73080 149336 73092
rect 123812 73052 149336 73080
rect 123812 73040 123818 73052
rect 149330 73040 149336 73052
rect 149388 73080 149394 73092
rect 149882 73080 149888 73092
rect 149388 73052 149888 73080
rect 149388 73040 149394 73052
rect 149882 73040 149888 73052
rect 149940 73040 149946 73092
rect 157518 73040 157524 73092
rect 157576 73080 157582 73092
rect 158530 73080 158536 73092
rect 157576 73052 158536 73080
rect 157576 73040 157582 73052
rect 158530 73040 158536 73052
rect 158588 73040 158594 73092
rect 165982 73040 165988 73092
rect 166040 73080 166046 73092
rect 198090 73080 198096 73092
rect 166040 73052 198096 73080
rect 166040 73040 166046 73052
rect 198090 73040 198096 73052
rect 198148 73080 198154 73092
rect 206278 73080 206284 73092
rect 198148 73052 206284 73080
rect 198148 73040 198154 73052
rect 206278 73040 206284 73052
rect 206336 73040 206342 73092
rect 119982 72972 119988 73024
rect 120040 73012 120046 73024
rect 151998 73012 152004 73024
rect 120040 72984 152004 73012
rect 120040 72972 120046 72984
rect 151998 72972 152004 72984
rect 152056 72972 152062 73024
rect 155678 72972 155684 73024
rect 155736 73012 155742 73024
rect 190086 73012 190092 73024
rect 155736 72984 190092 73012
rect 155736 72972 155742 72984
rect 190086 72972 190092 72984
rect 190144 72972 190150 73024
rect 106090 72904 106096 72956
rect 106148 72944 106154 72956
rect 139118 72944 139124 72956
rect 106148 72916 139124 72944
rect 106148 72904 106154 72916
rect 139118 72904 139124 72916
rect 139176 72904 139182 72956
rect 143994 72904 144000 72956
rect 144052 72944 144058 72956
rect 144270 72944 144276 72956
rect 144052 72916 144276 72944
rect 144052 72904 144058 72916
rect 144270 72904 144276 72916
rect 144328 72904 144334 72956
rect 163406 72904 163412 72956
rect 163464 72944 163470 72956
rect 163682 72944 163688 72956
rect 163464 72916 163688 72944
rect 163464 72904 163470 72916
rect 163682 72904 163688 72916
rect 163740 72904 163746 72956
rect 164694 72904 164700 72956
rect 164752 72944 164758 72956
rect 165430 72944 165436 72956
rect 164752 72916 165436 72944
rect 164752 72904 164758 72916
rect 165430 72904 165436 72916
rect 165488 72944 165494 72956
rect 199470 72944 199476 72956
rect 165488 72916 199476 72944
rect 165488 72904 165494 72916
rect 199470 72904 199476 72916
rect 199528 72904 199534 72956
rect 107470 72836 107476 72888
rect 107528 72876 107534 72888
rect 138566 72876 138572 72888
rect 107528 72848 138572 72876
rect 107528 72836 107534 72848
rect 138566 72836 138572 72848
rect 138624 72836 138630 72888
rect 155954 72836 155960 72888
rect 156012 72876 156018 72888
rect 156966 72876 156972 72888
rect 156012 72848 156972 72876
rect 156012 72836 156018 72848
rect 156966 72836 156972 72848
rect 157024 72836 157030 72888
rect 166994 72836 167000 72888
rect 167052 72876 167058 72888
rect 202414 72876 202420 72888
rect 167052 72848 202420 72876
rect 167052 72836 167058 72848
rect 202414 72836 202420 72848
rect 202472 72836 202478 72888
rect 111610 72768 111616 72820
rect 111668 72808 111674 72820
rect 143074 72808 143080 72820
rect 111668 72780 143080 72808
rect 111668 72768 111674 72780
rect 143074 72768 143080 72780
rect 143132 72768 143138 72820
rect 156598 72768 156604 72820
rect 156656 72808 156662 72820
rect 311158 72808 311164 72820
rect 156656 72780 311164 72808
rect 156656 72768 156662 72780
rect 311158 72768 311164 72780
rect 311216 72768 311222 72820
rect 104434 72700 104440 72752
rect 104492 72740 104498 72752
rect 130654 72740 130660 72752
rect 104492 72712 130660 72740
rect 104492 72700 104498 72712
rect 130654 72700 130660 72712
rect 130712 72700 130718 72752
rect 157242 72700 157248 72752
rect 157300 72740 157306 72752
rect 318794 72740 318800 72752
rect 157300 72712 318800 72740
rect 157300 72700 157306 72712
rect 318794 72700 318800 72712
rect 318852 72700 318858 72752
rect 115842 72632 115848 72684
rect 115900 72672 115906 72684
rect 141142 72672 141148 72684
rect 115900 72644 141148 72672
rect 115900 72632 115906 72644
rect 141142 72632 141148 72644
rect 141200 72632 141206 72684
rect 157702 72632 157708 72684
rect 157760 72672 157766 72684
rect 324958 72672 324964 72684
rect 157760 72644 324964 72672
rect 157760 72632 157766 72644
rect 324958 72632 324964 72644
rect 325016 72632 325022 72684
rect 70394 72564 70400 72616
rect 70452 72604 70458 72616
rect 137830 72604 137836 72616
rect 70452 72576 137836 72604
rect 70452 72564 70458 72576
rect 137830 72564 137836 72576
rect 137888 72564 137894 72616
rect 157610 72564 157616 72616
rect 157668 72604 157674 72616
rect 332594 72604 332600 72616
rect 157668 72576 332600 72604
rect 157668 72564 157674 72576
rect 332594 72564 332600 72576
rect 332652 72564 332658 72616
rect 23474 72496 23480 72548
rect 23532 72536 23538 72548
rect 100294 72536 100300 72548
rect 23532 72508 100300 72536
rect 23532 72496 23538 72508
rect 100294 72496 100300 72508
rect 100352 72536 100358 72548
rect 100352 72508 113174 72536
rect 100352 72496 100358 72508
rect 14458 72428 14464 72480
rect 14516 72468 14522 72480
rect 104434 72468 104440 72480
rect 14516 72440 104440 72468
rect 14516 72428 14522 72440
rect 104434 72428 104440 72440
rect 104492 72428 104498 72480
rect 113146 72264 113174 72508
rect 123938 72496 123944 72548
rect 123996 72536 124002 72548
rect 149514 72536 149520 72548
rect 123996 72508 149520 72536
rect 123996 72496 124002 72508
rect 149514 72496 149520 72508
rect 149572 72536 149578 72548
rect 149882 72536 149888 72548
rect 149572 72508 149888 72536
rect 149572 72496 149578 72508
rect 149882 72496 149888 72508
rect 149940 72496 149946 72548
rect 166166 72496 166172 72548
rect 166224 72536 166230 72548
rect 368474 72536 368480 72548
rect 166224 72508 368480 72536
rect 166224 72496 166230 72508
rect 368474 72496 368480 72508
rect 368532 72496 368538 72548
rect 116486 72428 116492 72480
rect 116544 72468 116550 72480
rect 141602 72468 141608 72480
rect 116544 72440 141608 72468
rect 116544 72428 116550 72440
rect 141602 72428 141608 72440
rect 141660 72428 141666 72480
rect 158254 72428 158260 72480
rect 158312 72468 158318 72480
rect 191098 72468 191104 72480
rect 158312 72440 191104 72468
rect 158312 72428 158318 72440
rect 191098 72428 191104 72440
rect 191156 72428 191162 72480
rect 202414 72428 202420 72480
rect 202472 72468 202478 72480
rect 446398 72468 446404 72480
rect 202472 72440 446404 72468
rect 202472 72428 202478 72440
rect 446398 72428 446404 72440
rect 446456 72428 446462 72480
rect 122742 72360 122748 72412
rect 122800 72400 122806 72412
rect 129918 72400 129924 72412
rect 122800 72372 129924 72400
rect 122800 72360 122806 72372
rect 129918 72360 129924 72372
rect 129976 72400 129982 72412
rect 132494 72400 132500 72412
rect 129976 72372 132500 72400
rect 129976 72360 129982 72372
rect 132494 72360 132500 72372
rect 132552 72360 132558 72412
rect 145006 72360 145012 72412
rect 145064 72400 145070 72412
rect 145374 72400 145380 72412
rect 145064 72372 145380 72400
rect 145064 72360 145070 72372
rect 145374 72360 145380 72372
rect 145432 72360 145438 72412
rect 158530 72360 158536 72412
rect 158588 72400 158594 72412
rect 189994 72400 190000 72412
rect 158588 72372 190000 72400
rect 158588 72360 158594 72372
rect 189994 72360 190000 72372
rect 190052 72360 190058 72412
rect 166994 72292 167000 72344
rect 167052 72332 167058 72344
rect 168098 72332 168104 72344
rect 167052 72304 168104 72332
rect 167052 72292 167058 72304
rect 168098 72292 168104 72304
rect 168156 72292 168162 72344
rect 176102 72292 176108 72344
rect 176160 72332 176166 72344
rect 204530 72332 204536 72344
rect 176160 72304 204536 72332
rect 176160 72292 176166 72304
rect 204530 72292 204536 72304
rect 204588 72292 204594 72344
rect 134334 72264 134340 72276
rect 113146 72236 134340 72264
rect 134334 72224 134340 72236
rect 134392 72224 134398 72276
rect 151998 72224 152004 72276
rect 152056 72264 152062 72276
rect 152826 72264 152832 72276
rect 152056 72236 152832 72264
rect 152056 72224 152062 72236
rect 152826 72224 152832 72236
rect 152884 72224 152890 72276
rect 161106 72224 161112 72276
rect 161164 72264 161170 72276
rect 187234 72264 187240 72276
rect 161164 72236 187240 72264
rect 161164 72224 161170 72236
rect 187234 72224 187240 72236
rect 187292 72224 187298 72276
rect 134334 72088 134340 72140
rect 134392 72128 134398 72140
rect 135162 72128 135168 72140
rect 134392 72100 135168 72128
rect 134392 72088 134398 72100
rect 135162 72088 135168 72100
rect 135220 72088 135226 72140
rect 175918 72088 175924 72140
rect 175976 72128 175982 72140
rect 176286 72128 176292 72140
rect 175976 72100 176292 72128
rect 175976 72088 175982 72100
rect 176286 72088 176292 72100
rect 176344 72088 176350 72140
rect 128906 71952 128912 72004
rect 128964 71992 128970 72004
rect 133230 71992 133236 72004
rect 128964 71964 133236 71992
rect 128964 71952 128970 71964
rect 133230 71952 133236 71964
rect 133288 71952 133294 72004
rect 115934 71748 115940 71800
rect 115992 71788 115998 71800
rect 116486 71788 116492 71800
rect 115992 71760 116492 71788
rect 115992 71748 115998 71760
rect 116486 71748 116492 71760
rect 116544 71748 116550 71800
rect 124950 71748 124956 71800
rect 125008 71788 125014 71800
rect 126238 71788 126244 71800
rect 125008 71760 126244 71788
rect 125008 71748 125014 71760
rect 126238 71748 126244 71760
rect 126296 71748 126302 71800
rect 127342 71748 127348 71800
rect 127400 71788 127406 71800
rect 127400 71760 127940 71788
rect 127400 71748 127406 71760
rect 122098 71680 122104 71732
rect 122156 71720 122162 71732
rect 122834 71720 122840 71732
rect 122156 71692 122840 71720
rect 122156 71680 122162 71692
rect 122834 71680 122840 71692
rect 122892 71680 122898 71732
rect 123294 71680 123300 71732
rect 123352 71720 123358 71732
rect 127434 71720 127440 71732
rect 123352 71692 127440 71720
rect 123352 71680 123358 71692
rect 127434 71680 127440 71692
rect 127492 71680 127498 71732
rect 127912 71720 127940 71760
rect 151906 71720 151912 71732
rect 127544 71692 127848 71720
rect 127912 71692 151912 71720
rect 3510 71612 3516 71664
rect 3568 71652 3574 71664
rect 8938 71652 8944 71664
rect 3568 71624 8944 71652
rect 3568 71612 3574 71624
rect 8938 71612 8944 71624
rect 8996 71612 9002 71664
rect 99374 71612 99380 71664
rect 99432 71652 99438 71664
rect 100386 71652 100392 71664
rect 99432 71624 100392 71652
rect 99432 71612 99438 71624
rect 100386 71612 100392 71624
rect 100444 71652 100450 71664
rect 127544 71652 127572 71692
rect 100444 71624 127572 71652
rect 127820 71652 127848 71692
rect 151906 71680 151912 71692
rect 151964 71680 151970 71732
rect 156414 71680 156420 71732
rect 156472 71720 156478 71732
rect 156690 71720 156696 71732
rect 156472 71692 156696 71720
rect 156472 71680 156478 71692
rect 156690 71680 156696 71692
rect 156748 71680 156754 71732
rect 159634 71680 159640 71732
rect 159692 71720 159698 71732
rect 160002 71720 160008 71732
rect 159692 71692 160008 71720
rect 159692 71680 159698 71692
rect 160002 71680 160008 71692
rect 160060 71680 160066 71732
rect 160830 71680 160836 71732
rect 160888 71720 160894 71732
rect 161290 71720 161296 71732
rect 160888 71692 161296 71720
rect 160888 71680 160894 71692
rect 161290 71680 161296 71692
rect 161348 71680 161354 71732
rect 161934 71680 161940 71732
rect 161992 71720 161998 71732
rect 162578 71720 162584 71732
rect 161992 71692 162584 71720
rect 161992 71680 161998 71692
rect 162578 71680 162584 71692
rect 162636 71680 162642 71732
rect 183646 71680 183652 71732
rect 183704 71720 183710 71732
rect 204438 71720 204444 71732
rect 183704 71692 204444 71720
rect 183704 71680 183710 71692
rect 204438 71680 204444 71692
rect 204496 71680 204502 71732
rect 134426 71652 134432 71664
rect 127820 71624 134432 71652
rect 100444 71612 100450 71624
rect 134426 71612 134432 71624
rect 134484 71612 134490 71664
rect 141418 71612 141424 71664
rect 141476 71652 141482 71664
rect 143074 71652 143080 71664
rect 141476 71624 143080 71652
rect 141476 71612 141482 71624
rect 143074 71612 143080 71624
rect 143132 71612 143138 71664
rect 151354 71612 151360 71664
rect 151412 71652 151418 71664
rect 151538 71652 151544 71664
rect 151412 71624 151544 71652
rect 151412 71612 151418 71624
rect 151538 71612 151544 71624
rect 151596 71612 151602 71664
rect 117498 71544 117504 71596
rect 117556 71584 117562 71596
rect 127342 71584 127348 71596
rect 117556 71556 127348 71584
rect 117556 71544 117562 71556
rect 127342 71544 127348 71556
rect 127400 71544 127406 71596
rect 127802 71544 127808 71596
rect 127860 71584 127866 71596
rect 156432 71584 156460 71680
rect 158806 71612 158812 71664
rect 158864 71652 158870 71664
rect 159726 71652 159732 71664
rect 158864 71624 159732 71652
rect 158864 71612 158870 71624
rect 159726 71612 159732 71624
rect 159784 71612 159790 71664
rect 160278 71612 160284 71664
rect 160336 71652 160342 71664
rect 161014 71652 161020 71664
rect 160336 71624 161020 71652
rect 160336 71612 160342 71624
rect 161014 71612 161020 71624
rect 161072 71652 161078 71664
rect 194962 71652 194968 71664
rect 161072 71624 194968 71652
rect 161072 71612 161078 71624
rect 194962 71612 194968 71624
rect 195020 71612 195026 71664
rect 127860 71556 156460 71584
rect 127860 71544 127866 71556
rect 162578 71544 162584 71596
rect 162636 71584 162642 71596
rect 196434 71584 196440 71596
rect 162636 71556 196440 71584
rect 162636 71544 162642 71556
rect 196434 71544 196440 71556
rect 196492 71544 196498 71596
rect 116946 71476 116952 71528
rect 117004 71516 117010 71528
rect 149790 71516 149796 71528
rect 117004 71488 149796 71516
rect 117004 71476 117010 71488
rect 149790 71476 149796 71488
rect 149848 71476 149854 71528
rect 158806 71476 158812 71528
rect 158864 71516 158870 71528
rect 159358 71516 159364 71528
rect 158864 71488 159364 71516
rect 158864 71476 158870 71488
rect 159358 71476 159364 71488
rect 159416 71476 159422 71528
rect 169662 71476 169668 71528
rect 169720 71516 169726 71528
rect 203518 71516 203524 71528
rect 169720 71488 203524 71516
rect 169720 71476 169726 71488
rect 203518 71476 203524 71488
rect 203576 71476 203582 71528
rect 108758 71408 108764 71460
rect 108816 71448 108822 71460
rect 140590 71448 140596 71460
rect 108816 71420 140596 71448
rect 108816 71408 108822 71420
rect 140590 71408 140596 71420
rect 140648 71408 140654 71460
rect 162118 71408 162124 71460
rect 162176 71448 162182 71460
rect 196894 71448 196900 71460
rect 162176 71420 196900 71448
rect 162176 71408 162182 71420
rect 196894 71408 196900 71420
rect 196952 71408 196958 71460
rect 120810 71340 120816 71392
rect 120868 71380 120874 71392
rect 152458 71380 152464 71392
rect 120868 71352 152464 71380
rect 120868 71340 120874 71352
rect 152458 71340 152464 71352
rect 152516 71340 152522 71392
rect 161290 71340 161296 71392
rect 161348 71380 161354 71392
rect 194226 71380 194232 71392
rect 161348 71352 194232 71380
rect 161348 71340 161354 71352
rect 194226 71340 194232 71352
rect 194284 71340 194290 71392
rect 119062 71272 119068 71324
rect 119120 71312 119126 71324
rect 119120 71284 147674 71312
rect 119120 71272 119126 71284
rect 120994 71204 121000 71256
rect 121052 71244 121058 71256
rect 147646 71244 147674 71284
rect 162394 71272 162400 71324
rect 162452 71312 162458 71324
rect 195422 71312 195428 71324
rect 162452 71284 195428 71312
rect 162452 71272 162458 71284
rect 195422 71272 195428 71284
rect 195480 71272 195486 71324
rect 151262 71244 151268 71256
rect 121052 71216 142844 71244
rect 147646 71216 151268 71244
rect 121052 71204 121058 71216
rect 27614 71136 27620 71188
rect 27672 71176 27678 71188
rect 99374 71176 99380 71188
rect 27672 71148 99380 71176
rect 27672 71136 27678 71148
rect 99374 71136 99380 71148
rect 99432 71136 99438 71188
rect 108942 71136 108948 71188
rect 109000 71176 109006 71188
rect 138198 71176 138204 71188
rect 109000 71148 138204 71176
rect 109000 71136 109006 71148
rect 138198 71136 138204 71148
rect 138256 71176 138262 71188
rect 139210 71176 139216 71188
rect 138256 71148 139216 71176
rect 138256 71136 138262 71148
rect 139210 71136 139216 71148
rect 139268 71136 139274 71188
rect 142816 71176 142844 71216
rect 151262 71204 151268 71216
rect 151320 71204 151326 71256
rect 159726 71204 159732 71256
rect 159784 71244 159790 71256
rect 192294 71244 192300 71256
rect 159784 71216 192300 71244
rect 159784 71204 159790 71216
rect 192294 71204 192300 71216
rect 192352 71204 192358 71256
rect 151354 71176 151360 71188
rect 142816 71148 151360 71176
rect 151354 71136 151360 71148
rect 151412 71136 151418 71188
rect 151906 71136 151912 71188
rect 151964 71176 151970 71188
rect 152642 71176 152648 71188
rect 151964 71148 152648 71176
rect 151964 71136 151970 71148
rect 152642 71136 152648 71148
rect 152700 71136 152706 71188
rect 166626 71136 166632 71188
rect 166684 71176 166690 71188
rect 166810 71176 166816 71188
rect 166684 71148 166816 71176
rect 166684 71136 166690 71148
rect 166810 71136 166816 71148
rect 166868 71176 166874 71188
rect 187142 71176 187148 71188
rect 166868 71148 187148 71176
rect 166868 71136 166874 71148
rect 187142 71136 187148 71148
rect 187200 71136 187206 71188
rect 26234 71068 26240 71120
rect 26292 71108 26298 71120
rect 102134 71108 102140 71120
rect 26292 71080 102140 71108
rect 26292 71068 26298 71080
rect 102134 71068 102140 71080
rect 102192 71068 102198 71120
rect 113450 71068 113456 71120
rect 113508 71108 113514 71120
rect 140406 71108 140412 71120
rect 113508 71080 140412 71108
rect 113508 71068 113514 71080
rect 140406 71068 140412 71080
rect 140464 71068 140470 71120
rect 148962 71068 148968 71120
rect 149020 71108 149026 71120
rect 179414 71108 179420 71120
rect 149020 71080 179420 71108
rect 149020 71068 149026 71080
rect 179414 71068 179420 71080
rect 179472 71068 179478 71120
rect 179506 71068 179512 71120
rect 179564 71108 179570 71120
rect 185026 71108 185032 71120
rect 179564 71080 185032 71108
rect 179564 71068 179570 71080
rect 185026 71068 185032 71080
rect 185084 71068 185090 71120
rect 185136 71080 186544 71108
rect 45554 71000 45560 71052
rect 45612 71040 45618 71052
rect 135990 71040 135996 71052
rect 45612 71012 135996 71040
rect 45612 71000 45618 71012
rect 135990 71000 135996 71012
rect 136048 71000 136054 71052
rect 160462 71000 160468 71052
rect 160520 71040 160526 71052
rect 185136 71040 185164 71080
rect 160520 71012 185164 71040
rect 186516 71040 186544 71080
rect 188338 71068 188344 71120
rect 188396 71108 188402 71120
rect 196618 71108 196624 71120
rect 188396 71080 196624 71108
rect 188396 71068 188402 71080
rect 196618 71068 196624 71080
rect 196676 71068 196682 71120
rect 204438 71068 204444 71120
rect 204496 71108 204502 71120
rect 218054 71108 218060 71120
rect 204496 71080 218060 71108
rect 204496 71068 204502 71080
rect 218054 71068 218060 71080
rect 218112 71068 218118 71120
rect 354674 71040 354680 71052
rect 186516 71012 354680 71040
rect 160520 71000 160526 71012
rect 354674 71000 354680 71012
rect 354732 71000 354738 71052
rect 117682 70932 117688 70984
rect 117740 70972 117746 70984
rect 136818 70972 136824 70984
rect 117740 70944 136824 70972
rect 117740 70932 117746 70944
rect 136818 70932 136824 70944
rect 136876 70972 136882 70984
rect 142890 70972 142896 70984
rect 136876 70944 142896 70972
rect 136876 70932 136882 70944
rect 142890 70932 142896 70944
rect 142948 70932 142954 70984
rect 160002 70932 160008 70984
rect 160060 70972 160066 70984
rect 160060 70944 166994 70972
rect 160060 70932 160066 70944
rect 114278 70864 114284 70916
rect 114336 70904 114342 70916
rect 128354 70904 128360 70916
rect 114336 70876 128360 70904
rect 114336 70864 114342 70876
rect 128354 70864 128360 70876
rect 128412 70904 128418 70916
rect 137094 70904 137100 70916
rect 128412 70876 137100 70904
rect 128412 70864 128418 70876
rect 137094 70864 137100 70876
rect 137152 70864 137158 70916
rect 160094 70864 160100 70916
rect 160152 70904 160158 70916
rect 160738 70904 160744 70916
rect 160152 70876 160744 70904
rect 160152 70864 160158 70876
rect 160738 70864 160744 70876
rect 160796 70864 160802 70916
rect 166966 70904 166994 70944
rect 180886 70932 180892 70984
rect 180944 70972 180950 70984
rect 188338 70972 188344 70984
rect 180944 70944 188344 70972
rect 180944 70932 180950 70944
rect 188338 70932 188344 70944
rect 188396 70932 188402 70984
rect 193950 70904 193956 70916
rect 166966 70876 193956 70904
rect 193950 70864 193956 70876
rect 194008 70864 194014 70916
rect 102134 70796 102140 70848
rect 102192 70836 102198 70848
rect 103054 70836 103060 70848
rect 102192 70808 103060 70836
rect 102192 70796 102198 70808
rect 103054 70796 103060 70808
rect 103112 70836 103118 70848
rect 129550 70836 129556 70848
rect 103112 70808 129556 70836
rect 103112 70796 103118 70808
rect 129550 70796 129556 70808
rect 129608 70796 129614 70848
rect 144270 70796 144276 70848
rect 144328 70836 144334 70848
rect 147122 70836 147128 70848
rect 144328 70808 147128 70836
rect 144328 70796 144334 70808
rect 147122 70796 147128 70808
rect 147180 70796 147186 70848
rect 189166 70728 189172 70780
rect 189224 70768 189230 70780
rect 189350 70768 189356 70780
rect 189224 70740 189356 70768
rect 189224 70728 189230 70740
rect 189350 70728 189356 70740
rect 189408 70728 189414 70780
rect 142522 70660 142528 70712
rect 142580 70700 142586 70712
rect 142982 70700 142988 70712
rect 142580 70672 142988 70700
rect 142580 70660 142586 70672
rect 142982 70660 142988 70672
rect 143040 70660 143046 70712
rect 107654 70388 107660 70440
rect 107712 70428 107718 70440
rect 108758 70428 108764 70440
rect 107712 70400 108764 70428
rect 107712 70388 107718 70400
rect 108758 70388 108764 70400
rect 108816 70388 108822 70440
rect 119614 70320 119620 70372
rect 119672 70360 119678 70372
rect 153194 70360 153200 70372
rect 119672 70332 153200 70360
rect 119672 70320 119678 70332
rect 153194 70320 153200 70332
rect 153252 70360 153258 70372
rect 153838 70360 153844 70372
rect 153252 70332 153844 70360
rect 153252 70320 153258 70332
rect 153838 70320 153844 70332
rect 153896 70320 153902 70372
rect 167178 70320 167184 70372
rect 167236 70360 167242 70372
rect 168098 70360 168104 70372
rect 167236 70332 168104 70360
rect 167236 70320 167242 70332
rect 168098 70320 168104 70332
rect 168156 70360 168162 70372
rect 202138 70360 202144 70372
rect 168156 70332 202144 70360
rect 168156 70320 168162 70332
rect 202138 70320 202144 70332
rect 202196 70320 202202 70372
rect 121730 70252 121736 70304
rect 121788 70292 121794 70304
rect 155218 70292 155224 70304
rect 121788 70264 155224 70292
rect 121788 70252 121794 70264
rect 155218 70252 155224 70264
rect 155276 70252 155282 70304
rect 167270 70252 167276 70304
rect 167328 70292 167334 70304
rect 167822 70292 167828 70304
rect 167328 70264 167828 70292
rect 167328 70252 167334 70264
rect 167822 70252 167828 70264
rect 167880 70292 167886 70304
rect 202230 70292 202236 70304
rect 167880 70264 202236 70292
rect 167880 70252 167886 70264
rect 202230 70252 202236 70264
rect 202288 70252 202294 70304
rect 120442 70184 120448 70236
rect 120500 70224 120506 70236
rect 153654 70224 153660 70236
rect 120500 70196 153660 70224
rect 120500 70184 120506 70196
rect 153654 70184 153660 70196
rect 153712 70224 153718 70236
rect 154206 70224 154212 70236
rect 153712 70196 154212 70224
rect 153712 70184 153718 70196
rect 154206 70184 154212 70196
rect 154264 70184 154270 70236
rect 162486 70184 162492 70236
rect 162544 70224 162550 70236
rect 196526 70224 196532 70236
rect 162544 70196 196532 70224
rect 162544 70184 162550 70196
rect 196526 70184 196532 70196
rect 196584 70184 196590 70236
rect 120902 70116 120908 70168
rect 120960 70156 120966 70168
rect 154114 70156 154120 70168
rect 120960 70128 154120 70156
rect 120960 70116 120966 70128
rect 154114 70116 154120 70128
rect 154172 70116 154178 70168
rect 164970 70116 164976 70168
rect 165028 70156 165034 70168
rect 199562 70156 199568 70168
rect 165028 70128 199568 70156
rect 165028 70116 165034 70128
rect 199562 70116 199568 70128
rect 199620 70116 199626 70168
rect 122006 70048 122012 70100
rect 122064 70088 122070 70100
rect 122064 70060 142154 70088
rect 122064 70048 122070 70060
rect 131574 70020 131580 70032
rect 103486 69992 131580 70020
rect 46198 69708 46204 69760
rect 46256 69748 46262 69760
rect 102962 69748 102968 69760
rect 46256 69720 102968 69748
rect 46256 69708 46262 69720
rect 102962 69708 102968 69720
rect 103020 69748 103026 69760
rect 103486 69748 103514 69992
rect 131574 69980 131580 69992
rect 131632 69980 131638 70032
rect 142126 70020 142154 70060
rect 144546 70048 144552 70100
rect 144604 70088 144610 70100
rect 146294 70088 146300 70100
rect 144604 70060 146300 70088
rect 144604 70048 144610 70060
rect 146294 70048 146300 70060
rect 146352 70048 146358 70100
rect 165338 70048 165344 70100
rect 165396 70088 165402 70100
rect 199654 70088 199660 70100
rect 165396 70060 199660 70088
rect 165396 70048 165402 70060
rect 199654 70048 199660 70060
rect 199712 70048 199718 70100
rect 153562 70020 153568 70032
rect 142126 69992 153568 70020
rect 153562 69980 153568 69992
rect 153620 70020 153626 70032
rect 153930 70020 153936 70032
rect 153620 69992 153936 70020
rect 153620 69980 153626 69992
rect 153930 69980 153936 69992
rect 153988 69980 153994 70032
rect 163866 69980 163872 70032
rect 163924 70020 163930 70032
rect 163924 69992 165108 70020
rect 163924 69980 163930 69992
rect 113542 69912 113548 69964
rect 113600 69952 113606 69964
rect 142522 69952 142528 69964
rect 113600 69924 142528 69952
rect 113600 69912 113606 69924
rect 142522 69912 142528 69924
rect 142580 69952 142586 69964
rect 143258 69952 143264 69964
rect 142580 69924 143264 69952
rect 142580 69912 142586 69924
rect 143258 69912 143264 69924
rect 143316 69912 143322 69964
rect 164326 69912 164332 69964
rect 164384 69952 164390 69964
rect 164970 69952 164976 69964
rect 164384 69924 164976 69952
rect 164384 69912 164390 69924
rect 164970 69912 164976 69924
rect 165028 69912 165034 69964
rect 165080 69952 165108 69992
rect 165154 69980 165160 70032
rect 165212 70020 165218 70032
rect 199378 70020 199384 70032
rect 165212 69992 199384 70020
rect 165212 69980 165218 69992
rect 199378 69980 199384 69992
rect 199436 69980 199442 70032
rect 198182 69952 198188 69964
rect 165080 69924 198188 69952
rect 198182 69912 198188 69924
rect 198240 69912 198246 69964
rect 112714 69844 112720 69896
rect 112772 69884 112778 69896
rect 139486 69884 139492 69896
rect 112772 69856 139492 69884
rect 112772 69844 112778 69856
rect 139486 69844 139492 69856
rect 139544 69844 139550 69896
rect 161658 69844 161664 69896
rect 161716 69884 161722 69896
rect 162486 69884 162492 69896
rect 161716 69856 162492 69884
rect 161716 69844 161722 69856
rect 162486 69844 162492 69856
rect 162544 69844 162550 69896
rect 164510 69844 164516 69896
rect 164568 69884 164574 69896
rect 165338 69884 165344 69896
rect 164568 69856 165344 69884
rect 164568 69844 164574 69856
rect 165338 69844 165344 69856
rect 165396 69844 165402 69896
rect 165890 69844 165896 69896
rect 165948 69884 165954 69896
rect 166626 69884 166632 69896
rect 165948 69856 166632 69884
rect 165948 69844 165954 69856
rect 166626 69844 166632 69856
rect 166684 69884 166690 69896
rect 200850 69884 200856 69896
rect 166684 69856 200856 69884
rect 166684 69844 166690 69856
rect 200850 69844 200856 69856
rect 200908 69844 200914 69896
rect 115014 69776 115020 69828
rect 115072 69816 115078 69828
rect 142154 69816 142160 69828
rect 115072 69788 142160 69816
rect 115072 69776 115078 69788
rect 142154 69776 142160 69788
rect 142212 69816 142218 69828
rect 142614 69816 142620 69828
rect 142212 69788 142620 69816
rect 142212 69776 142218 69788
rect 142614 69776 142620 69788
rect 142672 69776 142678 69828
rect 163038 69776 163044 69828
rect 163096 69816 163102 69828
rect 163866 69816 163872 69828
rect 163096 69788 163872 69816
rect 163096 69776 163102 69788
rect 163866 69776 163872 69788
rect 163924 69776 163930 69828
rect 164602 69776 164608 69828
rect 164660 69816 164666 69828
rect 165154 69816 165160 69828
rect 164660 69788 165160 69816
rect 164660 69776 164666 69788
rect 165154 69776 165160 69788
rect 165212 69776 165218 69828
rect 169110 69776 169116 69828
rect 169168 69816 169174 69828
rect 201770 69816 201776 69828
rect 169168 69788 201776 69816
rect 169168 69776 169174 69788
rect 201770 69776 201776 69788
rect 201828 69816 201834 69828
rect 202782 69816 202788 69828
rect 201828 69788 202788 69816
rect 201828 69776 201834 69788
rect 202782 69776 202788 69788
rect 202840 69776 202846 69828
rect 103020 69720 103514 69748
rect 103020 69708 103026 69720
rect 115566 69708 115572 69760
rect 115624 69748 115630 69760
rect 138106 69748 138112 69760
rect 115624 69720 138112 69748
rect 115624 69708 115630 69720
rect 138106 69708 138112 69720
rect 138164 69748 138170 69760
rect 138566 69748 138572 69760
rect 138164 69720 138572 69748
rect 138164 69708 138170 69720
rect 138566 69708 138572 69720
rect 138624 69708 138630 69760
rect 139486 69708 139492 69760
rect 139544 69748 139550 69760
rect 140314 69748 140320 69760
rect 139544 69720 140320 69748
rect 139544 69708 139550 69720
rect 140314 69708 140320 69720
rect 140372 69708 140378 69760
rect 164418 69708 164424 69760
rect 164476 69748 164482 69760
rect 188522 69748 188528 69760
rect 164476 69720 188528 69748
rect 164476 69708 164482 69720
rect 188522 69708 188528 69720
rect 188580 69748 188586 69760
rect 423766 69748 423772 69760
rect 188580 69720 423772 69748
rect 188580 69708 188586 69720
rect 423766 69708 423772 69720
rect 423824 69708 423830 69760
rect 18598 69640 18604 69692
rect 18656 69680 18662 69692
rect 18656 69652 84194 69680
rect 18656 69640 18662 69652
rect 84166 69612 84194 69652
rect 119798 69640 119804 69692
rect 119856 69680 119862 69692
rect 128446 69680 128452 69692
rect 119856 69652 128452 69680
rect 119856 69640 119862 69652
rect 128446 69640 128452 69652
rect 128504 69680 128510 69692
rect 142430 69680 142436 69692
rect 128504 69652 142436 69680
rect 128504 69640 128510 69652
rect 142430 69640 142436 69652
rect 142488 69640 142494 69692
rect 147950 69640 147956 69692
rect 148008 69680 148014 69692
rect 181530 69680 181536 69692
rect 148008 69652 181536 69680
rect 148008 69640 148014 69652
rect 181530 69640 181536 69652
rect 181588 69640 181594 69692
rect 202782 69640 202788 69692
rect 202840 69680 202846 69692
rect 448514 69680 448520 69692
rect 202840 69652 448520 69680
rect 202840 69640 202846 69652
rect 448514 69640 448520 69652
rect 448572 69640 448578 69692
rect 103146 69612 103152 69624
rect 84166 69584 103152 69612
rect 103146 69572 103152 69584
rect 103204 69612 103210 69624
rect 130194 69612 130200 69624
rect 103204 69584 130200 69612
rect 103204 69572 103210 69584
rect 130194 69572 130200 69584
rect 130252 69572 130258 69624
rect 103514 69504 103520 69556
rect 103572 69544 103578 69556
rect 108482 69544 108488 69556
rect 103572 69516 108488 69544
rect 103572 69504 103578 69516
rect 108482 69504 108488 69516
rect 108540 69504 108546 69556
rect 109034 68960 109040 69012
rect 109092 69000 109098 69012
rect 110966 69000 110972 69012
rect 109092 68972 110972 69000
rect 109092 68960 109098 68972
rect 110966 68960 110972 68972
rect 111024 68960 111030 69012
rect 118326 68960 118332 69012
rect 118384 69000 118390 69012
rect 152274 69000 152280 69012
rect 118384 68972 152280 69000
rect 118384 68960 118390 68972
rect 152274 68960 152280 68972
rect 152332 69000 152338 69012
rect 152550 69000 152556 69012
rect 152332 68972 152556 69000
rect 152332 68960 152338 68972
rect 152550 68960 152556 68972
rect 152608 68960 152614 69012
rect 167086 68960 167092 69012
rect 167144 69000 167150 69012
rect 168282 69000 168288 69012
rect 167144 68972 168288 69000
rect 167144 68960 167150 68972
rect 168282 68960 168288 68972
rect 168340 69000 168346 69012
rect 202046 69000 202052 69012
rect 168340 68972 202052 69000
rect 168340 68960 168346 68972
rect 202046 68960 202052 68972
rect 202104 68960 202110 69012
rect 117222 68892 117228 68944
rect 117280 68932 117286 68944
rect 151170 68932 151176 68944
rect 117280 68904 151176 68932
rect 117280 68892 117286 68904
rect 151170 68892 151176 68904
rect 151228 68892 151234 68944
rect 161474 68892 161480 68944
rect 161532 68932 161538 68944
rect 189166 68932 189172 68944
rect 161532 68904 189172 68932
rect 161532 68892 161538 68904
rect 189166 68892 189172 68904
rect 189224 68892 189230 68944
rect 108850 68824 108856 68876
rect 108908 68864 108914 68876
rect 142338 68864 142344 68876
rect 108908 68836 142344 68864
rect 108908 68824 108914 68836
rect 142338 68824 142344 68836
rect 142396 68864 142402 68876
rect 142706 68864 142712 68876
rect 142396 68836 142712 68864
rect 142396 68824 142402 68836
rect 142706 68824 142712 68836
rect 142764 68824 142770 68876
rect 176930 68824 176936 68876
rect 176988 68864 176994 68876
rect 199378 68864 199384 68876
rect 176988 68836 199384 68864
rect 176988 68824 176994 68836
rect 199378 68824 199384 68836
rect 199436 68824 199442 68876
rect 104618 68756 104624 68808
rect 104676 68796 104682 68808
rect 136082 68796 136088 68808
rect 104676 68768 136088 68796
rect 104676 68756 104682 68768
rect 136082 68756 136088 68768
rect 136140 68756 136146 68808
rect 163590 68756 163596 68808
rect 163648 68796 163654 68808
rect 183002 68796 183008 68808
rect 163648 68768 183008 68796
rect 163648 68756 163654 68768
rect 183002 68756 183008 68768
rect 183060 68796 183066 68808
rect 183462 68796 183468 68808
rect 183060 68768 183468 68796
rect 183060 68756 183066 68768
rect 183462 68756 183468 68768
rect 183520 68756 183526 68808
rect 89714 68552 89720 68604
rect 89772 68592 89778 68604
rect 105722 68592 105728 68604
rect 89772 68564 105728 68592
rect 89772 68552 89778 68564
rect 105722 68552 105728 68564
rect 105780 68552 105786 68604
rect 131022 68552 131028 68604
rect 131080 68592 131086 68604
rect 135254 68592 135260 68604
rect 131080 68564 135260 68592
rect 131080 68552 131086 68564
rect 135254 68552 135260 68564
rect 135312 68552 135318 68604
rect 85574 68484 85580 68536
rect 85632 68524 85638 68536
rect 106090 68524 106096 68536
rect 85632 68496 106096 68524
rect 85632 68484 85638 68496
rect 106090 68484 106096 68496
rect 106148 68484 106154 68536
rect 120074 68484 120080 68536
rect 120132 68524 120138 68536
rect 141786 68524 141792 68536
rect 120132 68496 141792 68524
rect 120132 68484 120138 68496
rect 141786 68484 141792 68496
rect 141844 68484 141850 68536
rect 78674 68416 78680 68468
rect 78732 68456 78738 68468
rect 107470 68456 107476 68468
rect 78732 68428 107476 68456
rect 78732 68416 78738 68428
rect 107470 68416 107476 68428
rect 107528 68416 107534 68468
rect 118602 68416 118608 68468
rect 118660 68456 118666 68468
rect 141234 68456 141240 68468
rect 118660 68428 141240 68456
rect 118660 68416 118666 68428
rect 141234 68416 141240 68428
rect 141292 68416 141298 68468
rect 149882 68416 149888 68468
rect 149940 68456 149946 68468
rect 220814 68456 220820 68468
rect 149940 68428 220820 68456
rect 149940 68416 149946 68428
rect 220814 68416 220820 68428
rect 220872 68416 220878 68468
rect 75914 68348 75920 68400
rect 75972 68388 75978 68400
rect 107010 68388 107016 68400
rect 75972 68360 107016 68388
rect 75972 68348 75978 68360
rect 107010 68348 107016 68360
rect 107068 68348 107074 68400
rect 117314 68348 117320 68400
rect 117372 68388 117378 68400
rect 140958 68388 140964 68400
rect 117372 68360 140964 68388
rect 117372 68348 117378 68360
rect 140958 68348 140964 68360
rect 141016 68348 141022 68400
rect 189166 68348 189172 68400
rect 189224 68388 189230 68400
rect 302234 68388 302240 68400
rect 189224 68360 302240 68388
rect 189224 68348 189230 68360
rect 302234 68348 302240 68360
rect 302292 68348 302298 68400
rect 48314 68280 48320 68332
rect 48372 68320 48378 68332
rect 104618 68320 104624 68332
rect 48372 68292 104624 68320
rect 48372 68280 48378 68292
rect 104618 68280 104624 68292
rect 104676 68280 104682 68332
rect 113174 68280 113180 68332
rect 113232 68320 113238 68332
rect 140774 68320 140780 68332
rect 113232 68292 140780 68320
rect 113232 68280 113238 68292
rect 140774 68280 140780 68292
rect 140832 68280 140838 68332
rect 186682 68280 186688 68332
rect 186740 68320 186746 68332
rect 504358 68320 504364 68332
rect 186740 68292 504364 68320
rect 186740 68280 186746 68292
rect 504358 68280 504364 68292
rect 504416 68280 504422 68332
rect 183462 67668 183468 67720
rect 183520 67708 183526 67720
rect 332686 67708 332692 67720
rect 183520 67680 332692 67708
rect 183520 67668 183526 67680
rect 332686 67668 332692 67680
rect 332744 67668 332750 67720
rect 199378 67600 199384 67652
rect 199436 67640 199442 67652
rect 560938 67640 560944 67652
rect 199436 67612 560944 67640
rect 199436 67600 199442 67612
rect 560938 67600 560944 67612
rect 560996 67600 561002 67652
rect 104342 67532 104348 67584
rect 104400 67572 104406 67584
rect 138474 67572 138480 67584
rect 104400 67544 138480 67572
rect 104400 67532 104406 67544
rect 138474 67532 138480 67544
rect 138532 67532 138538 67584
rect 144914 67532 144920 67584
rect 144972 67572 144978 67584
rect 147214 67572 147220 67584
rect 144972 67544 147220 67572
rect 144972 67532 144978 67544
rect 147214 67532 147220 67544
rect 147272 67532 147278 67584
rect 165798 67532 165804 67584
rect 165856 67572 165862 67584
rect 200390 67572 200396 67584
rect 165856 67544 200396 67572
rect 165856 67532 165862 67544
rect 200390 67532 200396 67544
rect 200448 67572 200454 67584
rect 201402 67572 201408 67584
rect 200448 67544 201408 67572
rect 200448 67532 200454 67544
rect 201402 67532 201408 67544
rect 201460 67532 201466 67584
rect 114002 67464 114008 67516
rect 114060 67504 114066 67516
rect 139854 67504 139860 67516
rect 114060 67476 139860 67504
rect 114060 67464 114066 67476
rect 139854 67464 139860 67476
rect 139912 67464 139918 67516
rect 110138 67396 110144 67448
rect 110196 67436 110202 67448
rect 118602 67436 118608 67448
rect 110196 67408 118608 67436
rect 110196 67396 110202 67408
rect 118602 67396 118608 67408
rect 118660 67396 118666 67448
rect 92474 67124 92480 67176
rect 92532 67164 92538 67176
rect 105630 67164 105636 67176
rect 92532 67136 105636 67164
rect 92532 67124 92538 67136
rect 105630 67124 105636 67136
rect 105688 67124 105694 67176
rect 93946 67056 93952 67108
rect 94004 67096 94010 67108
rect 112530 67096 112536 67108
rect 94004 67068 112536 67096
rect 94004 67056 94010 67068
rect 112530 67056 112536 67068
rect 112588 67056 112594 67108
rect 80054 66988 80060 67040
rect 80112 67028 80118 67040
rect 104342 67028 104348 67040
rect 80112 67000 104348 67028
rect 80112 66988 80118 67000
rect 104342 66988 104348 67000
rect 104400 66988 104406 67040
rect 106274 66988 106280 67040
rect 106332 67028 106338 67040
rect 139578 67028 139584 67040
rect 106332 67000 139584 67028
rect 106332 66988 106338 67000
rect 139578 66988 139584 67000
rect 139636 66988 139642 67040
rect 102134 66920 102140 66972
rect 102192 66960 102198 66972
rect 139670 66960 139676 66972
rect 102192 66932 139676 66960
rect 102192 66920 102198 66932
rect 139670 66920 139676 66932
rect 139728 66920 139734 66972
rect 164786 66920 164792 66972
rect 164844 66960 164850 66972
rect 389174 66960 389180 66972
rect 164844 66932 389180 66960
rect 164844 66920 164850 66932
rect 389174 66920 389180 66932
rect 389232 66920 389238 66972
rect 99374 66852 99380 66904
rect 99432 66892 99438 66904
rect 139762 66892 139768 66904
rect 99432 66864 139768 66892
rect 99432 66852 99438 66864
rect 139762 66852 139768 66864
rect 139820 66852 139826 66904
rect 201402 66852 201408 66904
rect 201460 66892 201466 66904
rect 432598 66892 432604 66904
rect 201460 66864 432604 66892
rect 201460 66852 201466 66864
rect 432598 66852 432604 66864
rect 432656 66852 432662 66904
rect 140774 66240 140780 66292
rect 140832 66280 140838 66292
rect 142154 66280 142160 66292
rect 140832 66252 142160 66280
rect 140832 66240 140838 66252
rect 142154 66240 142160 66252
rect 142212 66240 142218 66292
rect 189166 66240 189172 66292
rect 189224 66280 189230 66292
rect 539594 66280 539600 66292
rect 189224 66252 539600 66280
rect 189224 66240 189230 66252
rect 539594 66240 539600 66252
rect 539652 66240 539658 66292
rect 102226 66172 102232 66224
rect 102284 66212 102290 66224
rect 103238 66212 103244 66224
rect 102284 66184 103244 66212
rect 102284 66172 102290 66184
rect 103238 66172 103244 66184
rect 103296 66212 103302 66224
rect 134334 66212 134340 66224
rect 103296 66184 134340 66212
rect 103296 66172 103302 66184
rect 134334 66172 134340 66184
rect 134392 66172 134398 66224
rect 143994 66172 144000 66224
rect 144052 66212 144058 66224
rect 148410 66212 148416 66224
rect 144052 66184 148416 66212
rect 144052 66172 144058 66184
rect 148410 66172 148416 66184
rect 148468 66172 148474 66224
rect 159082 66172 159088 66224
rect 159140 66212 159146 66224
rect 190914 66212 190920 66224
rect 159140 66184 190920 66212
rect 159140 66172 159146 66184
rect 190914 66172 190920 66184
rect 190972 66212 190978 66224
rect 191742 66212 191748 66224
rect 190972 66184 191748 66212
rect 190972 66172 190978 66184
rect 191742 66172 191748 66184
rect 191800 66172 191806 66224
rect 97994 65560 98000 65612
rect 98052 65600 98058 65612
rect 111058 65600 111064 65612
rect 98052 65572 111064 65600
rect 98052 65560 98058 65572
rect 111058 65560 111064 65572
rect 111116 65560 111122 65612
rect 148778 65560 148784 65612
rect 148836 65600 148842 65612
rect 207014 65600 207020 65612
rect 148836 65572 207020 65600
rect 148836 65560 148842 65572
rect 207014 65560 207020 65572
rect 207072 65560 207078 65612
rect 35986 65492 35992 65544
rect 36044 65532 36050 65544
rect 102226 65532 102232 65544
rect 36044 65504 102232 65532
rect 36044 65492 36050 65504
rect 102226 65492 102232 65504
rect 102284 65492 102290 65544
rect 146478 65492 146484 65544
rect 146536 65532 146542 65544
rect 183554 65532 183560 65544
rect 146536 65504 183560 65532
rect 146536 65492 146542 65504
rect 183554 65492 183560 65504
rect 183612 65492 183618 65544
rect 191742 65492 191748 65544
rect 191800 65532 191806 65544
rect 346394 65532 346400 65544
rect 191800 65504 346400 65532
rect 191800 65492 191806 65504
rect 346394 65492 346400 65504
rect 346452 65492 346458 65544
rect 139394 64880 139400 64932
rect 139452 64920 139458 64932
rect 142154 64920 142160 64932
rect 139452 64892 142160 64920
rect 139452 64880 139458 64892
rect 142154 64880 142160 64892
rect 142212 64880 142218 64932
rect 102226 64812 102232 64864
rect 102284 64852 102290 64864
rect 103330 64852 103336 64864
rect 102284 64824 103336 64852
rect 102284 64812 102290 64824
rect 103330 64812 103336 64824
rect 103388 64852 103394 64864
rect 137186 64852 137192 64864
rect 103388 64824 137192 64852
rect 103388 64812 103394 64824
rect 137186 64812 137192 64824
rect 137244 64812 137250 64864
rect 168834 64812 168840 64864
rect 168892 64852 168898 64864
rect 203058 64852 203064 64864
rect 168892 64824 203064 64852
rect 168892 64812 168898 64824
rect 203058 64812 203064 64824
rect 203116 64812 203122 64864
rect 149698 64268 149704 64320
rect 149756 64308 149762 64320
rect 224954 64308 224960 64320
rect 149756 64280 224960 64308
rect 149756 64268 149762 64280
rect 224954 64268 224960 64280
rect 225012 64268 225018 64320
rect 62114 64200 62120 64252
rect 62172 64240 62178 64252
rect 102226 64240 102232 64252
rect 62172 64212 102232 64240
rect 62172 64200 62178 64212
rect 102226 64200 102232 64212
rect 102284 64200 102290 64252
rect 152826 64200 152832 64252
rect 152884 64240 152890 64252
rect 256694 64240 256700 64252
rect 152884 64212 256700 64240
rect 152884 64200 152890 64212
rect 256694 64200 256700 64212
rect 256752 64200 256758 64252
rect 4154 64132 4160 64184
rect 4212 64172 4218 64184
rect 132494 64172 132500 64184
rect 4212 64144 132500 64172
rect 4212 64132 4218 64144
rect 132494 64132 132500 64144
rect 132552 64132 132558 64184
rect 150526 64132 150532 64184
rect 150584 64172 150590 64184
rect 183002 64172 183008 64184
rect 150584 64144 183008 64172
rect 150584 64132 150590 64144
rect 183002 64132 183008 64144
rect 183060 64132 183066 64184
rect 203058 64132 203064 64184
rect 203116 64172 203122 64184
rect 472618 64172 472624 64184
rect 203116 64144 472624 64172
rect 203116 64132 203122 64144
rect 472618 64132 472624 64144
rect 472676 64132 472682 64184
rect 104710 63452 104716 63504
rect 104768 63492 104774 63504
rect 132770 63492 132776 63504
rect 104768 63464 132776 63492
rect 104768 63452 104774 63464
rect 132770 63452 132776 63464
rect 132828 63452 132834 63504
rect 158990 63452 158996 63504
rect 159048 63492 159054 63504
rect 193214 63492 193220 63504
rect 159048 63464 193220 63492
rect 159048 63452 159054 63464
rect 193214 63452 193220 63464
rect 193272 63452 193278 63504
rect 88334 62840 88340 62892
rect 88392 62880 88398 62892
rect 138382 62880 138388 62892
rect 88392 62852 138388 62880
rect 88392 62840 88398 62852
rect 138382 62840 138388 62852
rect 138440 62840 138446 62892
rect 193214 62840 193220 62892
rect 193272 62880 193278 62892
rect 340874 62880 340880 62892
rect 193272 62852 340880 62880
rect 193272 62840 193278 62852
rect 340874 62840 340880 62852
rect 340932 62840 340938 62892
rect 10318 62772 10324 62824
rect 10376 62812 10382 62824
rect 104710 62812 104716 62824
rect 10376 62784 104716 62812
rect 10376 62772 10382 62784
rect 104710 62772 104716 62784
rect 104768 62772 104774 62824
rect 160186 62772 160192 62824
rect 160244 62812 160250 62824
rect 357434 62812 357440 62824
rect 160244 62784 357440 62812
rect 160244 62772 160250 62784
rect 357434 62772 357440 62784
rect 357492 62772 357498 62824
rect 102226 62024 102232 62076
rect 102284 62064 102290 62076
rect 103422 62064 103428 62076
rect 102284 62036 103428 62064
rect 102284 62024 102290 62036
rect 103422 62024 103428 62036
rect 103480 62064 103486 62076
rect 135806 62064 135812 62076
rect 103480 62036 135812 62064
rect 103480 62024 103486 62036
rect 135806 62024 135812 62036
rect 135864 62024 135870 62076
rect 162946 62024 162952 62076
rect 163004 62064 163010 62076
rect 197354 62064 197360 62076
rect 163004 62036 197360 62064
rect 163004 62024 163010 62036
rect 197354 62024 197360 62036
rect 197412 62064 197418 62076
rect 197538 62064 197544 62076
rect 197412 62036 197544 62064
rect 197412 62024 197418 62036
rect 197538 62024 197544 62036
rect 197596 62024 197602 62076
rect 166350 61956 166356 62008
rect 166408 61996 166414 62008
rect 197630 61996 197636 62008
rect 166408 61968 197636 61996
rect 166408 61956 166414 61968
rect 197630 61956 197636 61968
rect 197688 61956 197694 62008
rect 135346 61888 135352 61940
rect 135404 61928 135410 61940
rect 142982 61928 142988 61940
rect 135404 61900 142988 61928
rect 135404 61888 135410 61900
rect 142982 61888 142988 61900
rect 143040 61888 143046 61940
rect 176838 61888 176844 61940
rect 176896 61928 176902 61940
rect 196066 61928 196072 61940
rect 176896 61900 196072 61928
rect 176896 61888 176902 61900
rect 196066 61888 196072 61900
rect 196124 61888 196130 61940
rect 172698 61820 172704 61872
rect 172756 61860 172762 61872
rect 186958 61860 186964 61872
rect 172756 61832 186964 61860
rect 172756 61820 172762 61832
rect 186958 61820 186964 61832
rect 187016 61820 187022 61872
rect 144638 61480 144644 61532
rect 144696 61520 144702 61532
rect 149698 61520 149704 61532
rect 144696 61492 149704 61520
rect 144696 61480 144702 61492
rect 149698 61480 149704 61492
rect 149756 61480 149762 61532
rect 52546 61412 52552 61464
rect 52604 61452 52610 61464
rect 102226 61452 102232 61464
rect 52604 61424 102232 61452
rect 52604 61412 52610 61424
rect 102226 61412 102232 61424
rect 102284 61412 102290 61464
rect 197354 61412 197360 61464
rect 197412 61452 197418 61464
rect 394694 61452 394700 61464
rect 197412 61424 394700 61452
rect 197412 61412 197418 61424
rect 394694 61412 394700 61424
rect 394752 61412 394758 61464
rect 42794 61344 42800 61396
rect 42852 61384 42858 61396
rect 135714 61384 135720 61396
rect 42852 61356 135720 61384
rect 42852 61344 42858 61356
rect 135714 61344 135720 61356
rect 135772 61344 135778 61396
rect 197630 61344 197636 61396
rect 197688 61384 197694 61396
rect 198366 61384 198372 61396
rect 197688 61356 198372 61384
rect 197688 61344 197694 61356
rect 198366 61344 198372 61356
rect 198424 61384 198430 61396
rect 396074 61384 396080 61396
rect 198424 61356 396080 61384
rect 198424 61344 198430 61356
rect 396074 61344 396080 61356
rect 396132 61344 396138 61396
rect 186958 60800 186964 60852
rect 187016 60840 187022 60852
rect 529934 60840 529940 60852
rect 187016 60812 529940 60840
rect 187016 60800 187022 60812
rect 529934 60800 529940 60812
rect 529992 60800 529998 60852
rect 196066 60732 196072 60784
rect 196124 60772 196130 60784
rect 574738 60772 574744 60784
rect 196124 60744 574744 60772
rect 196124 60732 196130 60744
rect 574738 60732 574744 60744
rect 574796 60732 574802 60784
rect 99466 60664 99472 60716
rect 99524 60704 99530 60716
rect 100570 60704 100576 60716
rect 99524 60676 100576 60704
rect 99524 60664 99530 60676
rect 100570 60664 100576 60676
rect 100628 60704 100634 60716
rect 133598 60704 133604 60716
rect 100628 60676 133604 60704
rect 100628 60664 100634 60676
rect 133598 60664 133604 60676
rect 133656 60664 133662 60716
rect 158898 60664 158904 60716
rect 158956 60704 158962 60716
rect 193306 60704 193312 60716
rect 158956 60676 193312 60704
rect 158956 60664 158962 60676
rect 193306 60664 193312 60676
rect 193364 60704 193370 60716
rect 194502 60704 194508 60716
rect 193364 60676 194508 60704
rect 193364 60664 193370 60676
rect 194502 60664 194508 60676
rect 194560 60664 194566 60716
rect 104802 60596 104808 60648
rect 104860 60636 104866 60648
rect 137462 60636 137468 60648
rect 104860 60608 137468 60636
rect 104860 60596 104866 60608
rect 137462 60596 137468 60608
rect 137520 60596 137526 60648
rect 149790 60188 149796 60240
rect 149848 60228 149854 60240
rect 223574 60228 223580 60240
rect 149848 60200 223580 60228
rect 149848 60188 149854 60200
rect 223574 60188 223580 60200
rect 223632 60188 223638 60240
rect 145190 60120 145196 60172
rect 145248 60160 145254 60172
rect 147306 60160 147312 60172
rect 145248 60132 147312 60160
rect 145248 60120 145254 60132
rect 147306 60120 147312 60132
rect 147364 60120 147370 60172
rect 150802 60120 150808 60172
rect 150860 60160 150866 60172
rect 245654 60160 245660 60172
rect 150860 60132 245660 60160
rect 150860 60120 150866 60132
rect 245654 60120 245660 60132
rect 245712 60120 245718 60172
rect 69014 60052 69020 60104
rect 69072 60092 69078 60104
rect 104802 60092 104808 60104
rect 69072 60064 104808 60092
rect 69072 60052 69078 60064
rect 104802 60052 104808 60064
rect 104860 60052 104866 60104
rect 155310 60052 155316 60104
rect 155368 60092 155374 60104
rect 299474 60092 299480 60104
rect 155368 60064 299480 60092
rect 155368 60052 155374 60064
rect 299474 60052 299480 60064
rect 299532 60052 299538 60104
rect 17954 59984 17960 60036
rect 18012 60024 18018 60036
rect 99466 60024 99472 60036
rect 18012 59996 99472 60024
rect 18012 59984 18018 59996
rect 99466 59984 99472 59996
rect 99524 59984 99530 60036
rect 153102 59984 153108 60036
rect 153160 60024 153166 60036
rect 186314 60024 186320 60036
rect 153160 59996 186320 60024
rect 153160 59984 153166 59996
rect 186314 59984 186320 59996
rect 186372 59984 186378 60036
rect 194502 59984 194508 60036
rect 194560 60024 194566 60036
rect 345014 60024 345020 60036
rect 194560 59996 345020 60024
rect 194560 59984 194566 59996
rect 345014 59984 345020 59996
rect 345072 59984 345078 60036
rect 110414 59304 110420 59356
rect 110472 59344 110478 59356
rect 115198 59344 115204 59356
rect 110472 59316 115204 59344
rect 110472 59304 110478 59316
rect 115198 59304 115204 59316
rect 115256 59304 115262 59356
rect 135990 59344 135996 59356
rect 122806 59316 135996 59344
rect 111794 59236 111800 59288
rect 111852 59276 111858 59288
rect 112254 59276 112260 59288
rect 111852 59248 112260 59276
rect 111852 59236 111858 59248
rect 112254 59236 112260 59248
rect 112312 59276 112318 59288
rect 122806 59276 122834 59316
rect 135990 59304 135996 59316
rect 136048 59304 136054 59356
rect 112312 59248 122834 59276
rect 112312 59236 112318 59248
rect 147398 58692 147404 58744
rect 147456 58732 147462 58744
rect 193306 58732 193312 58744
rect 147456 58704 193312 58732
rect 147456 58692 147462 58704
rect 193306 58692 193312 58704
rect 193364 58692 193370 58744
rect 49694 58624 49700 58676
rect 49752 58664 49758 58676
rect 111794 58664 111800 58676
rect 49752 58636 111800 58664
rect 49752 58624 49758 58636
rect 111794 58624 111800 58636
rect 111852 58624 111858 58676
rect 170490 58624 170496 58676
rect 170548 58664 170554 58676
rect 490006 58664 490012 58676
rect 170548 58636 490012 58664
rect 170548 58624 170554 58636
rect 490006 58624 490012 58636
rect 490064 58624 490070 58676
rect 168742 57876 168748 57928
rect 168800 57916 168806 57928
rect 203426 57916 203432 57928
rect 168800 57888 203432 57916
rect 168800 57876 168806 57888
rect 203426 57876 203432 57888
rect 203484 57916 203490 57928
rect 204162 57916 204168 57928
rect 203484 57888 204168 57916
rect 203484 57876 203490 57888
rect 204162 57876 204168 57888
rect 204220 57876 204226 57928
rect 151446 57264 151452 57316
rect 151504 57304 151510 57316
rect 233234 57304 233240 57316
rect 151504 57276 233240 57304
rect 151504 57264 151510 57276
rect 233234 57264 233240 57276
rect 233292 57264 233298 57316
rect 204162 57196 204168 57248
rect 204220 57236 204226 57248
rect 473446 57236 473452 57248
rect 204220 57208 473452 57236
rect 204220 57196 204226 57208
rect 473446 57196 473452 57208
rect 473504 57196 473510 57248
rect 99466 56516 99472 56568
rect 99524 56556 99530 56568
rect 100662 56556 100668 56568
rect 99524 56528 100668 56556
rect 99524 56516 99530 56528
rect 100662 56516 100668 56528
rect 100720 56556 100726 56568
rect 133414 56556 133420 56568
rect 100720 56528 133420 56556
rect 100720 56516 100726 56528
rect 133414 56516 133420 56528
rect 133472 56516 133478 56568
rect 63494 55904 63500 55956
rect 63552 55944 63558 55956
rect 137002 55944 137008 55956
rect 63552 55916 137008 55944
rect 63552 55904 63558 55916
rect 137002 55904 137008 55916
rect 137060 55904 137066 55956
rect 147858 55904 147864 55956
rect 147916 55944 147922 55956
rect 197354 55944 197360 55956
rect 147916 55916 197360 55944
rect 147916 55904 147922 55916
rect 197354 55904 197360 55916
rect 197412 55904 197418 55956
rect 12434 55836 12440 55888
rect 12492 55876 12498 55888
rect 99466 55876 99472 55888
rect 12492 55848 99472 55876
rect 12492 55836 12498 55848
rect 99466 55836 99472 55848
rect 99524 55836 99530 55888
rect 148686 55836 148692 55888
rect 148744 55876 148750 55888
rect 204254 55876 204260 55888
rect 148744 55848 204260 55876
rect 148744 55836 148750 55848
rect 204254 55836 204260 55848
rect 204312 55836 204318 55888
rect 138658 55224 138664 55276
rect 138716 55264 138722 55276
rect 142338 55264 142344 55276
rect 138716 55236 142344 55264
rect 138716 55224 138722 55236
rect 142338 55224 142344 55236
rect 142396 55224 142402 55276
rect 168650 55156 168656 55208
rect 168708 55196 168714 55208
rect 201678 55196 201684 55208
rect 168708 55168 201684 55196
rect 168708 55156 168714 55168
rect 201678 55156 201684 55168
rect 201736 55196 201742 55208
rect 202782 55196 202788 55208
rect 201736 55168 202788 55196
rect 201736 55156 201742 55168
rect 202782 55156 202788 55168
rect 202840 55156 202846 55208
rect 148134 54544 148140 54596
rect 148192 54584 148198 54596
rect 209866 54584 209872 54596
rect 148192 54556 209872 54584
rect 148192 54544 148198 54556
rect 209866 54544 209872 54556
rect 209924 54544 209930 54596
rect 171042 54476 171048 54528
rect 171100 54516 171106 54528
rect 486418 54516 486424 54528
rect 171100 54488 486424 54516
rect 171100 54476 171106 54488
rect 486418 54476 486424 54488
rect 486476 54476 486482 54528
rect 202782 53796 202788 53848
rect 202840 53836 202846 53848
rect 464338 53836 464344 53848
rect 202840 53808 464344 53836
rect 202840 53796 202846 53808
rect 464338 53796 464344 53808
rect 464396 53796 464402 53848
rect 100478 53728 100484 53780
rect 100536 53768 100542 53780
rect 133046 53768 133052 53780
rect 100536 53740 133052 53768
rect 100536 53728 100542 53740
rect 133046 53728 133052 53740
rect 133104 53728 133110 53780
rect 168558 53728 168564 53780
rect 168616 53768 168622 53780
rect 203794 53768 203800 53780
rect 168616 53740 203800 53768
rect 168616 53728 168622 53740
rect 203794 53728 203800 53740
rect 203852 53728 203858 53780
rect 149238 53184 149244 53236
rect 149296 53224 149302 53236
rect 215294 53224 215300 53236
rect 149296 53196 215300 53224
rect 149296 53184 149302 53196
rect 215294 53184 215300 53196
rect 215352 53184 215358 53236
rect 157978 53116 157984 53168
rect 158036 53156 158042 53168
rect 333974 53156 333980 53168
rect 158036 53128 333980 53156
rect 158036 53116 158042 53128
rect 333974 53116 333980 53128
rect 334032 53116 334038 53168
rect 9674 53048 9680 53100
rect 9732 53088 9738 53100
rect 100478 53088 100484 53100
rect 9732 53060 100484 53088
rect 9732 53048 9738 53060
rect 100478 53048 100484 53060
rect 100536 53048 100542 53100
rect 102226 53048 102232 53100
rect 102284 53088 102290 53100
rect 113818 53088 113824 53100
rect 102284 53060 113824 53088
rect 102284 53048 102290 53060
rect 113818 53048 113824 53060
rect 113876 53048 113882 53100
rect 203794 53048 203800 53100
rect 203852 53088 203858 53100
rect 466454 53088 466460 53100
rect 203852 53060 466460 53088
rect 203852 53048 203858 53060
rect 466454 53048 466460 53060
rect 466512 53048 466518 53100
rect 169202 52368 169208 52420
rect 169260 52408 169266 52420
rect 202966 52408 202972 52420
rect 169260 52380 202972 52408
rect 169260 52368 169266 52380
rect 202966 52368 202972 52380
rect 203024 52408 203030 52420
rect 204162 52408 204168 52420
rect 203024 52380 204168 52408
rect 203024 52368 203030 52380
rect 204162 52368 204168 52380
rect 204220 52368 204226 52420
rect 145098 51824 145104 51876
rect 145156 51864 145162 51876
rect 169018 51864 169024 51876
rect 145156 51836 169024 51864
rect 145156 51824 145162 51836
rect 169018 51824 169024 51836
rect 169076 51824 169082 51876
rect 155954 51756 155960 51808
rect 156012 51796 156018 51808
rect 320174 51796 320180 51808
rect 156012 51768 320180 51796
rect 156012 51756 156018 51768
rect 320174 51756 320180 51768
rect 320232 51756 320238 51808
rect 147582 51688 147588 51740
rect 147640 51728 147646 51740
rect 191834 51728 191840 51740
rect 147640 51700 191840 51728
rect 147640 51688 147646 51700
rect 191834 51688 191840 51700
rect 191892 51688 191898 51740
rect 204162 51688 204168 51740
rect 204220 51728 204226 51740
rect 468478 51728 468484 51740
rect 204220 51700 468484 51728
rect 204220 51688 204226 51700
rect 468478 51688 468484 51700
rect 468536 51688 468542 51740
rect 100754 51008 100760 51060
rect 100812 51048 100818 51060
rect 105538 51048 105544 51060
rect 100812 51020 105544 51048
rect 100812 51008 100818 51020
rect 105538 51008 105544 51020
rect 105596 51008 105602 51060
rect 176746 51008 176752 51060
rect 176804 51048 176810 51060
rect 203058 51048 203064 51060
rect 176804 51020 203064 51048
rect 176804 51008 176810 51020
rect 203058 51008 203064 51020
rect 203116 51048 203122 51060
rect 204162 51048 204168 51060
rect 203116 51020 204168 51048
rect 203116 51008 203122 51020
rect 204162 51008 204168 51020
rect 204220 51008 204226 51060
rect 150158 50464 150164 50516
rect 150216 50504 150222 50516
rect 218146 50504 218152 50516
rect 150216 50476 218152 50504
rect 150216 50464 150222 50476
rect 218146 50464 218152 50476
rect 218204 50464 218210 50516
rect 152734 50396 152740 50448
rect 152792 50436 152798 50448
rect 259454 50436 259460 50448
rect 152792 50408 259460 50436
rect 152792 50396 152798 50408
rect 259454 50396 259460 50408
rect 259512 50396 259518 50448
rect 176654 50328 176660 50380
rect 176712 50368 176718 50380
rect 578234 50368 578240 50380
rect 176712 50340 578240 50368
rect 176712 50328 176718 50340
rect 578234 50328 578240 50340
rect 578292 50328 578298 50380
rect 204162 49716 204168 49768
rect 204220 49756 204226 49768
rect 569954 49756 569960 49768
rect 204220 49728 569960 49756
rect 204220 49716 204226 49728
rect 569954 49716 569960 49728
rect 570012 49716 570018 49768
rect 150250 49104 150256 49156
rect 150308 49144 150314 49156
rect 222194 49144 222200 49156
rect 150308 49116 222200 49144
rect 150308 49104 150314 49116
rect 222194 49104 222200 49116
rect 222252 49104 222258 49156
rect 155218 49036 155224 49088
rect 155276 49076 155282 49088
rect 285674 49076 285680 49088
rect 155276 49048 285680 49076
rect 155276 49036 155282 49048
rect 285674 49036 285680 49048
rect 285732 49036 285738 49088
rect 175274 48968 175280 49020
rect 175332 49008 175338 49020
rect 556154 49008 556160 49020
rect 175332 48980 556160 49008
rect 175332 48968 175338 48980
rect 556154 48968 556160 48980
rect 556212 48968 556218 49020
rect 147766 47744 147772 47796
rect 147824 47784 147830 47796
rect 201586 47784 201592 47796
rect 147824 47756 201592 47784
rect 147824 47744 147830 47756
rect 201586 47744 201592 47756
rect 201644 47744 201650 47796
rect 148594 47676 148600 47728
rect 148652 47716 148658 47728
rect 208394 47716 208400 47728
rect 148652 47688 208400 47716
rect 148652 47676 148658 47688
rect 208394 47676 208400 47688
rect 208452 47676 208458 47728
rect 170582 47608 170588 47660
rect 170640 47648 170646 47660
rect 488534 47648 488540 47660
rect 170640 47620 488540 47648
rect 170640 47608 170646 47620
rect 488534 47608 488540 47620
rect 488592 47608 488598 47660
rect 145006 47540 145012 47592
rect 145064 47580 145070 47592
rect 168558 47580 168564 47592
rect 145064 47552 168564 47580
rect 145064 47540 145070 47552
rect 168558 47540 168564 47552
rect 168616 47540 168622 47592
rect 177666 47540 177672 47592
rect 177724 47580 177730 47592
rect 582374 47580 582380 47592
rect 177724 47552 582380 47580
rect 177724 47540 177730 47552
rect 582374 47540 582380 47552
rect 582432 47540 582438 47592
rect 143810 46860 143816 46912
rect 143868 46900 143874 46912
rect 147766 46900 147772 46912
rect 143868 46872 147772 46900
rect 143868 46860 143874 46872
rect 147766 46860 147772 46872
rect 147824 46860 147830 46912
rect 177482 46860 177488 46912
rect 177540 46900 177546 46912
rect 204346 46900 204352 46912
rect 177540 46872 204352 46900
rect 177540 46860 177546 46872
rect 204346 46860 204352 46872
rect 204404 46900 204410 46912
rect 204714 46900 204720 46912
rect 204404 46872 204720 46900
rect 204404 46860 204410 46872
rect 204714 46860 204720 46872
rect 204772 46860 204778 46912
rect 151354 46384 151360 46436
rect 151412 46424 151418 46436
rect 235994 46424 236000 46436
rect 151412 46396 236000 46424
rect 151412 46384 151418 46396
rect 235994 46384 236000 46396
rect 236052 46384 236058 46436
rect 154298 46316 154304 46368
rect 154356 46356 154362 46368
rect 275278 46356 275284 46368
rect 154356 46328 275284 46356
rect 154356 46316 154362 46328
rect 275278 46316 275284 46328
rect 275336 46316 275342 46368
rect 168374 46248 168380 46300
rect 168432 46288 168438 46300
rect 474734 46288 474740 46300
rect 168432 46260 474740 46288
rect 168432 46248 168438 46260
rect 474734 46248 474740 46260
rect 474792 46248 474798 46300
rect 204714 46180 204720 46232
rect 204772 46220 204778 46232
rect 571978 46220 571984 46232
rect 204772 46192 571984 46220
rect 204772 46180 204778 46192
rect 571978 46180 571984 46192
rect 572036 46180 572042 46232
rect 161566 44956 161572 45008
rect 161624 44996 161630 45008
rect 390554 44996 390560 45008
rect 161624 44968 390560 44996
rect 161624 44956 161630 44968
rect 390554 44956 390560 44968
rect 390612 44956 390618 45008
rect 172514 44888 172520 44940
rect 172572 44928 172578 44940
rect 527174 44928 527180 44940
rect 172572 44900 527180 44928
rect 172572 44888 172578 44900
rect 527174 44888 527180 44900
rect 527232 44888 527238 44940
rect 60826 44820 60832 44872
rect 60884 44860 60890 44872
rect 137922 44860 137928 44872
rect 60884 44832 137928 44860
rect 60884 44820 60890 44832
rect 137922 44820 137928 44832
rect 137980 44820 137986 44872
rect 174630 44820 174636 44872
rect 174688 44860 174694 44872
rect 542354 44860 542360 44872
rect 174688 44832 542360 44860
rect 174688 44820 174694 44832
rect 542354 44820 542360 44832
rect 542412 44820 542418 44872
rect 156322 43528 156328 43580
rect 156380 43568 156386 43580
rect 315298 43568 315304 43580
rect 156380 43540 315304 43568
rect 156380 43528 156386 43540
rect 315298 43528 315304 43540
rect 315356 43528 315362 43580
rect 163774 43460 163780 43512
rect 163832 43500 163838 43512
rect 404354 43500 404360 43512
rect 163832 43472 404360 43500
rect 163832 43460 163838 43472
rect 404354 43460 404360 43472
rect 404412 43460 404418 43512
rect 162854 43392 162860 43444
rect 162912 43432 162918 43444
rect 408494 43432 408500 43444
rect 162912 43404 408500 43432
rect 162912 43392 162918 43404
rect 408494 43392 408500 43404
rect 408552 43392 408558 43444
rect 138014 42576 138020 42628
rect 138072 42616 138078 42628
rect 142246 42616 142252 42628
rect 138072 42588 142252 42616
rect 138072 42576 138078 42588
rect 142246 42576 142252 42588
rect 142304 42576 142310 42628
rect 155402 42304 155408 42356
rect 155460 42344 155466 42356
rect 292666 42344 292672 42356
rect 155460 42316 292672 42344
rect 155460 42304 155466 42316
rect 292666 42304 292672 42316
rect 292724 42304 292730 42356
rect 164234 42236 164240 42288
rect 164292 42276 164298 42288
rect 426434 42276 426440 42288
rect 164292 42248 426440 42276
rect 164292 42236 164298 42248
rect 426434 42236 426440 42248
rect 426492 42236 426498 42288
rect 166534 42168 166540 42220
rect 166592 42208 166598 42220
rect 440326 42208 440332 42220
rect 166592 42180 440332 42208
rect 166592 42168 166598 42180
rect 440326 42168 440332 42180
rect 440384 42168 440390 42220
rect 171318 42100 171324 42152
rect 171376 42140 171382 42152
rect 498286 42140 498292 42152
rect 171376 42112 498292 42140
rect 171376 42100 171382 42112
rect 498286 42100 498292 42112
rect 498344 42100 498350 42152
rect 77386 42032 77392 42084
rect 77444 42072 77450 42084
rect 138842 42072 138848 42084
rect 77444 42044 138848 42072
rect 77444 42032 77450 42044
rect 138842 42032 138848 42044
rect 138900 42032 138906 42084
rect 173618 42032 173624 42084
rect 173676 42072 173682 42084
rect 528554 42072 528560 42084
rect 173676 42044 528560 42072
rect 173676 42032 173682 42044
rect 528554 42032 528560 42044
rect 528612 42032 528618 42084
rect 148502 40944 148508 40996
rect 148560 40984 148566 40996
rect 205634 40984 205640 40996
rect 148560 40956 205640 40984
rect 148560 40944 148566 40956
rect 205634 40944 205640 40956
rect 205692 40944 205698 40996
rect 157058 40876 157064 40928
rect 157116 40916 157122 40928
rect 317414 40916 317420 40928
rect 157116 40888 317420 40916
rect 157116 40876 157122 40888
rect 317414 40876 317420 40888
rect 317472 40876 317478 40928
rect 165706 40808 165712 40860
rect 165764 40848 165770 40860
rect 444374 40848 444380 40860
rect 165764 40820 444380 40848
rect 165764 40808 165770 40820
rect 444374 40808 444380 40820
rect 444432 40808 444438 40860
rect 173434 40740 173440 40792
rect 173492 40780 173498 40792
rect 516134 40780 516140 40792
rect 173492 40752 516140 40780
rect 173492 40740 173498 40752
rect 516134 40740 516140 40752
rect 516192 40740 516198 40792
rect 13814 40672 13820 40724
rect 13872 40712 13878 40724
rect 132862 40712 132868 40724
rect 13872 40684 132868 40712
rect 13872 40672 13878 40684
rect 132862 40672 132868 40684
rect 132920 40672 132926 40724
rect 176194 40672 176200 40724
rect 176252 40712 176258 40724
rect 564526 40712 564532 40724
rect 176252 40684 564532 40712
rect 176252 40672 176258 40684
rect 564526 40672 564532 40684
rect 564584 40672 564590 40724
rect 152642 39584 152648 39636
rect 152700 39624 152706 39636
rect 251174 39624 251180 39636
rect 152700 39596 251180 39624
rect 152700 39584 152706 39596
rect 251174 39584 251180 39596
rect 251232 39584 251238 39636
rect 160738 39516 160744 39568
rect 160796 39556 160802 39568
rect 361574 39556 361580 39568
rect 160796 39528 361580 39556
rect 160796 39516 160802 39528
rect 361574 39516 361580 39528
rect 361632 39516 361638 39568
rect 168466 39448 168472 39500
rect 168524 39488 168530 39500
rect 463694 39488 463700 39500
rect 168524 39460 463700 39488
rect 168524 39448 168530 39460
rect 463694 39448 463700 39460
rect 463752 39448 463758 39500
rect 166994 39380 167000 39432
rect 167052 39420 167058 39432
rect 462314 39420 462320 39432
rect 167052 39392 462320 39420
rect 167052 39380 167058 39392
rect 462314 39380 462320 39392
rect 462372 39380 462378 39432
rect 31754 39312 31760 39364
rect 31812 39352 31818 39364
rect 134242 39352 134248 39364
rect 31812 39324 134248 39352
rect 31812 39312 31818 39324
rect 134242 39312 134248 39324
rect 134300 39312 134306 39364
rect 173526 39312 173532 39364
rect 173584 39352 173590 39364
rect 520274 39352 520280 39364
rect 173584 39324 520280 39352
rect 173584 39312 173590 39324
rect 520274 39312 520280 39324
rect 520332 39312 520338 39364
rect 154666 38156 154672 38208
rect 154724 38196 154730 38208
rect 293954 38196 293960 38208
rect 154724 38168 293960 38196
rect 154724 38156 154730 38168
rect 293954 38156 293960 38168
rect 294012 38156 294018 38208
rect 158806 38088 158812 38140
rect 158864 38128 158870 38140
rect 351914 38128 351920 38140
rect 158864 38100 351920 38128
rect 158864 38088 158870 38100
rect 351914 38088 351920 38100
rect 351972 38088 351978 38140
rect 167822 38020 167828 38072
rect 167880 38060 167886 38072
rect 448606 38060 448612 38072
rect 167880 38032 448612 38060
rect 167880 38020 167886 38032
rect 448606 38020 448612 38032
rect 448664 38020 448670 38072
rect 170674 37952 170680 38004
rect 170732 37992 170738 38004
rect 481634 37992 481640 38004
rect 170732 37964 481640 37992
rect 170732 37952 170738 37964
rect 481634 37952 481640 37964
rect 481692 37952 481698 38004
rect 38654 37884 38660 37936
rect 38712 37924 38718 37936
rect 135622 37924 135628 37936
rect 38712 37896 135628 37924
rect 38712 37884 38718 37896
rect 135622 37884 135628 37896
rect 135680 37884 135686 37936
rect 143718 37884 143724 37936
rect 143776 37924 143782 37936
rect 154574 37924 154580 37936
rect 143776 37896 154580 37924
rect 143776 37884 143782 37896
rect 154574 37884 154580 37896
rect 154632 37884 154638 37936
rect 174722 37884 174728 37936
rect 174780 37924 174786 37936
rect 538214 37924 538220 37936
rect 174780 37896 538220 37924
rect 174780 37884 174786 37896
rect 538214 37884 538220 37896
rect 538272 37884 538278 37936
rect 149054 36728 149060 36780
rect 149112 36768 149118 36780
rect 226334 36768 226340 36780
rect 149112 36740 226340 36768
rect 149112 36728 149118 36740
rect 226334 36728 226340 36740
rect 226392 36728 226398 36780
rect 155494 36660 155500 36712
rect 155552 36700 155558 36712
rect 299566 36700 299572 36712
rect 155552 36672 299572 36700
rect 155552 36660 155558 36672
rect 299566 36660 299572 36672
rect 299624 36660 299630 36712
rect 170766 36592 170772 36644
rect 170824 36632 170830 36644
rect 484394 36632 484400 36644
rect 170824 36604 484400 36632
rect 170824 36592 170830 36604
rect 484394 36592 484400 36604
rect 484452 36592 484458 36644
rect 176102 36524 176108 36576
rect 176160 36564 176166 36576
rect 552014 36564 552020 36576
rect 176160 36536 552020 36564
rect 176160 36524 176166 36536
rect 552014 36524 552020 36536
rect 552072 36524 552078 36576
rect 156874 35436 156880 35488
rect 156932 35476 156938 35488
rect 310514 35476 310520 35488
rect 156932 35448 310520 35476
rect 156932 35436 156938 35448
rect 310514 35436 310520 35448
rect 310572 35436 310578 35488
rect 159726 35368 159732 35420
rect 159784 35408 159790 35420
rect 342254 35408 342260 35420
rect 159784 35380 342260 35408
rect 159784 35368 159790 35380
rect 342254 35368 342260 35380
rect 342312 35368 342318 35420
rect 167914 35300 167920 35352
rect 167972 35340 167978 35352
rect 454034 35340 454040 35352
rect 167972 35312 454040 35340
rect 167972 35300 167978 35312
rect 454034 35300 454040 35312
rect 454092 35300 454098 35352
rect 171778 35232 171784 35284
rect 171836 35272 171842 35284
rect 502334 35272 502340 35284
rect 171836 35244 502340 35272
rect 171836 35232 171842 35244
rect 502334 35232 502340 35244
rect 502392 35232 502398 35284
rect 53834 35164 53840 35216
rect 53892 35204 53898 35216
rect 135438 35204 135444 35216
rect 53892 35176 135444 35204
rect 53892 35164 53898 35176
rect 135438 35164 135444 35176
rect 135496 35164 135502 35216
rect 144914 35164 144920 35216
rect 144972 35204 144978 35216
rect 166994 35204 167000 35216
rect 144972 35176 167000 35204
rect 144972 35164 144978 35176
rect 166994 35164 167000 35176
rect 167052 35164 167058 35216
rect 177758 35164 177764 35216
rect 177816 35204 177822 35216
rect 571334 35204 571340 35216
rect 177816 35176 571340 35204
rect 177816 35164 177822 35176
rect 571334 35164 571340 35176
rect 571392 35164 571398 35216
rect 152550 34008 152556 34060
rect 152608 34048 152614 34060
rect 251266 34048 251272 34060
rect 152608 34020 251272 34048
rect 152608 34008 152614 34020
rect 251266 34008 251272 34020
rect 251324 34008 251330 34060
rect 163866 33940 163872 33992
rect 163924 33980 163930 33992
rect 391934 33980 391940 33992
rect 163924 33952 391940 33980
rect 163924 33940 163930 33952
rect 391934 33940 391940 33952
rect 391992 33940 391998 33992
rect 165062 33872 165068 33924
rect 165120 33912 165126 33924
rect 410518 33912 410524 33924
rect 165120 33884 410524 33912
rect 165120 33872 165126 33884
rect 410518 33872 410524 33884
rect 410576 33872 410582 33924
rect 170858 33804 170864 33856
rect 170916 33844 170922 33856
rect 491294 33844 491300 33856
rect 170916 33816 491300 33844
rect 170916 33804 170922 33816
rect 491294 33804 491300 33816
rect 491352 33804 491358 33856
rect 177850 33736 177856 33788
rect 177908 33776 177914 33788
rect 576854 33776 576860 33788
rect 177908 33748 576860 33776
rect 177908 33736 177914 33748
rect 576854 33736 576860 33748
rect 576912 33736 576918 33788
rect 178954 33056 178960 33108
rect 179012 33096 179018 33108
rect 580166 33096 580172 33108
rect 179012 33068 580172 33096
rect 179012 33056 179018 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 154206 32580 154212 32632
rect 154264 32620 154270 32632
rect 267826 32620 267832 32632
rect 154264 32592 267832 32620
rect 154264 32580 154270 32592
rect 267826 32580 267832 32592
rect 267884 32580 267890 32632
rect 161014 32512 161020 32564
rect 161072 32552 161078 32564
rect 357526 32552 357532 32564
rect 161072 32524 357532 32552
rect 161072 32512 161078 32524
rect 357526 32512 357532 32524
rect 357584 32512 357590 32564
rect 166718 32444 166724 32496
rect 166776 32484 166782 32496
rect 431954 32484 431960 32496
rect 166776 32456 431960 32484
rect 166776 32444 166782 32456
rect 431954 32444 431960 32456
rect 432012 32444 432018 32496
rect 174814 32376 174820 32428
rect 174872 32416 174878 32428
rect 539686 32416 539692 32428
rect 174872 32388 539692 32416
rect 174872 32376 174878 32388
rect 539686 32376 539692 32388
rect 539744 32376 539750 32428
rect 148870 31356 148876 31408
rect 148928 31396 148934 31408
rect 198734 31396 198740 31408
rect 148928 31368 198740 31396
rect 148928 31356 148934 31368
rect 198734 31356 198740 31368
rect 198792 31356 198798 31408
rect 157150 31288 157156 31340
rect 157208 31328 157214 31340
rect 303614 31328 303620 31340
rect 157208 31300 303620 31328
rect 157208 31288 157214 31300
rect 303614 31288 303620 31300
rect 303672 31288 303678 31340
rect 163682 31220 163688 31272
rect 163740 31260 163746 31272
rect 340966 31260 340972 31272
rect 163740 31232 340972 31260
rect 163740 31220 163746 31232
rect 340966 31220 340972 31232
rect 341024 31220 341030 31272
rect 164970 31152 164976 31204
rect 165028 31192 165034 31204
rect 409874 31192 409880 31204
rect 165028 31164 409880 31192
rect 165028 31152 165034 31164
rect 409874 31152 409880 31164
rect 409932 31152 409938 31204
rect 183094 31084 183100 31136
rect 183152 31124 183158 31136
rect 442994 31124 443000 31136
rect 183152 31096 443000 31124
rect 183152 31084 183158 31096
rect 442994 31084 443000 31096
rect 443052 31084 443058 31136
rect 44266 31016 44272 31068
rect 44324 31056 44330 31068
rect 135530 31056 135536 31068
rect 44324 31028 135536 31056
rect 44324 31016 44330 31028
rect 135530 31016 135536 31028
rect 135588 31016 135594 31068
rect 169846 31016 169852 31068
rect 169904 31056 169910 31068
rect 495434 31056 495440 31068
rect 169904 31028 495440 31056
rect 169904 31016 169910 31028
rect 495434 31016 495440 31028
rect 495492 31016 495498 31068
rect 158254 29860 158260 29912
rect 158312 29900 158318 29912
rect 321554 29900 321560 29912
rect 158312 29872 321560 29900
rect 158312 29860 158318 29872
rect 321554 29860 321560 29872
rect 321612 29860 321618 29912
rect 167730 29792 167736 29844
rect 167788 29832 167794 29844
rect 375374 29832 375380 29844
rect 167788 29804 375380 29832
rect 167788 29792 167794 29804
rect 375374 29792 375380 29804
rect 375432 29792 375438 29844
rect 166626 29724 166632 29776
rect 166684 29764 166690 29776
rect 434714 29764 434720 29776
rect 166684 29736 434720 29764
rect 166684 29724 166690 29736
rect 434714 29724 434720 29736
rect 434772 29724 434778 29776
rect 177298 29656 177304 29708
rect 177356 29696 177362 29708
rect 554774 29696 554780 29708
rect 177356 29668 554780 29696
rect 177356 29656 177362 29668
rect 554774 29656 554780 29668
rect 554832 29656 554838 29708
rect 175366 29588 175372 29640
rect 175424 29628 175430 29640
rect 558178 29628 558184 29640
rect 175424 29600 558184 29628
rect 175424 29588 175430 29600
rect 558178 29588 558184 29600
rect 558236 29588 558242 29640
rect 143626 28908 143632 28960
rect 143684 28948 143690 28960
rect 144914 28948 144920 28960
rect 143684 28920 144920 28948
rect 143684 28908 143690 28920
rect 144914 28908 144920 28920
rect 144972 28908 144978 28960
rect 151262 28500 151268 28552
rect 151320 28540 151326 28552
rect 242986 28540 242992 28552
rect 151320 28512 242992 28540
rect 151320 28500 151326 28512
rect 242986 28500 242992 28512
rect 243044 28500 243050 28552
rect 159818 28432 159824 28484
rect 159876 28472 159882 28484
rect 339494 28472 339500 28484
rect 159876 28444 339500 28472
rect 159876 28432 159882 28444
rect 339494 28432 339500 28444
rect 339552 28432 339558 28484
rect 162026 28364 162032 28416
rect 162084 28404 162090 28416
rect 379514 28404 379520 28416
rect 162084 28376 379520 28404
rect 162084 28364 162090 28376
rect 379514 28364 379520 28376
rect 379572 28364 379578 28416
rect 168006 28296 168012 28348
rect 168064 28336 168070 28348
rect 456886 28336 456892 28348
rect 168064 28308 456892 28336
rect 168064 28296 168070 28308
rect 456886 28296 456892 28308
rect 456944 28296 456950 28348
rect 171962 28228 171968 28280
rect 172020 28268 172026 28280
rect 506566 28268 506572 28280
rect 172020 28240 506572 28268
rect 172020 28228 172026 28240
rect 506566 28228 506572 28240
rect 506624 28228 506630 28280
rect 162302 27072 162308 27124
rect 162360 27112 162366 27124
rect 374086 27112 374092 27124
rect 162360 27084 374092 27112
rect 162360 27072 162366 27084
rect 374086 27072 374092 27084
rect 374144 27072 374150 27124
rect 178862 27004 178868 27056
rect 178920 27044 178926 27056
rect 407114 27044 407120 27056
rect 178920 27016 407120 27044
rect 178920 27004 178926 27016
rect 407114 27004 407120 27016
rect 407172 27004 407178 27056
rect 172146 26936 172152 26988
rect 172204 26976 172210 26988
rect 509234 26976 509240 26988
rect 172204 26948 509240 26976
rect 172204 26936 172210 26948
rect 509234 26936 509240 26948
rect 509292 26936 509298 26988
rect 173710 26868 173716 26920
rect 173768 26908 173774 26920
rect 524414 26908 524420 26920
rect 173768 26880 524420 26908
rect 173768 26868 173774 26880
rect 524414 26868 524420 26880
rect 524472 26868 524478 26920
rect 154022 25780 154028 25832
rect 154080 25820 154086 25832
rect 278774 25820 278780 25832
rect 154080 25792 278780 25820
rect 154080 25780 154086 25792
rect 278774 25780 278780 25792
rect 278832 25780 278838 25832
rect 162394 25712 162400 25764
rect 162452 25752 162458 25764
rect 382366 25752 382372 25764
rect 162452 25724 382372 25752
rect 162452 25712 162458 25724
rect 382366 25712 382372 25724
rect 382424 25712 382430 25764
rect 165246 25644 165252 25696
rect 165304 25684 165310 25696
rect 425054 25684 425060 25696
rect 165304 25656 425060 25684
rect 165304 25644 165310 25656
rect 425054 25644 425060 25656
rect 425112 25644 425118 25696
rect 172238 25576 172244 25628
rect 172296 25616 172302 25628
rect 513374 25616 513380 25628
rect 172296 25588 513380 25616
rect 172296 25576 172302 25588
rect 513374 25576 513380 25588
rect 513432 25576 513438 25628
rect 173250 25508 173256 25560
rect 173308 25548 173314 25560
rect 531406 25548 531412 25560
rect 173308 25520 531412 25548
rect 173308 25508 173314 25520
rect 531406 25508 531412 25520
rect 531464 25508 531470 25560
rect 154114 24284 154120 24336
rect 154172 24324 154178 24336
rect 282914 24324 282920 24336
rect 154172 24296 282920 24324
rect 154172 24284 154178 24296
rect 282914 24284 282920 24296
rect 282972 24284 282978 24336
rect 163958 24216 163964 24268
rect 164016 24256 164022 24268
rect 398926 24256 398932 24268
rect 164016 24228 398932 24256
rect 164016 24216 164022 24228
rect 398926 24216 398932 24228
rect 398984 24216 398990 24268
rect 173158 24148 173164 24200
rect 173216 24188 173222 24200
rect 522298 24188 522304 24200
rect 173216 24160 522304 24188
rect 173216 24148 173222 24160
rect 522298 24148 522304 24160
rect 522356 24148 522362 24200
rect 146202 24080 146208 24132
rect 146260 24120 146266 24132
rect 173250 24120 173256 24132
rect 146260 24092 173256 24120
rect 146260 24080 146266 24092
rect 173250 24080 173256 24092
rect 173308 24080 173314 24132
rect 174998 24080 175004 24132
rect 175056 24120 175062 24132
rect 546494 24120 546500 24132
rect 175056 24092 546500 24120
rect 175056 24080 175062 24092
rect 546494 24080 546500 24092
rect 546552 24080 546558 24132
rect 149974 22992 149980 23044
rect 150032 23032 150038 23044
rect 219434 23032 219440 23044
rect 150032 23004 219440 23032
rect 150032 22992 150038 23004
rect 219434 22992 219440 23004
rect 219492 22992 219498 23044
rect 159910 22924 159916 22976
rect 159968 22964 159974 22976
rect 350534 22964 350540 22976
rect 159968 22936 350540 22964
rect 159968 22924 159974 22936
rect 350534 22924 350540 22936
rect 350592 22924 350598 22976
rect 165154 22856 165160 22908
rect 165212 22896 165218 22908
rect 416774 22896 416780 22908
rect 165212 22868 416780 22896
rect 165212 22856 165218 22868
rect 416774 22856 416780 22868
rect 416832 22856 416838 22908
rect 168190 22788 168196 22840
rect 168248 22828 168254 22840
rect 460934 22828 460940 22840
rect 168248 22800 460940 22828
rect 168248 22788 168254 22800
rect 460934 22788 460940 22800
rect 460992 22788 460998 22840
rect 174906 22720 174912 22772
rect 174964 22760 174970 22772
rect 534074 22760 534080 22772
rect 174964 22732 534080 22760
rect 174964 22720 174970 22732
rect 534074 22720 534080 22732
rect 534132 22720 534138 22772
rect 157794 21564 157800 21616
rect 157852 21604 157858 21616
rect 322934 21604 322940 21616
rect 157852 21576 322940 21604
rect 157852 21564 157858 21576
rect 322934 21564 322940 21576
rect 322992 21564 322998 21616
rect 158346 21496 158352 21548
rect 158404 21536 158410 21548
rect 329834 21536 329840 21548
rect 158404 21508 329840 21536
rect 158404 21496 158410 21508
rect 329834 21496 329840 21508
rect 329892 21496 329898 21548
rect 158438 21428 158444 21480
rect 158496 21468 158502 21480
rect 336734 21468 336740 21480
rect 158496 21440 336740 21468
rect 158496 21428 158502 21440
rect 336734 21428 336740 21440
rect 336792 21428 336798 21480
rect 337378 21428 337384 21480
rect 337436 21468 337442 21480
rect 471974 21468 471980 21480
rect 337436 21440 471980 21468
rect 337436 21428 337442 21440
rect 471974 21428 471980 21440
rect 472032 21428 472038 21480
rect 158714 21360 158720 21412
rect 158772 21400 158778 21412
rect 343634 21400 343640 21412
rect 158772 21372 343640 21400
rect 158772 21360 158778 21372
rect 343634 21360 343640 21372
rect 343692 21360 343698 21412
rect 289078 20612 289084 20664
rect 289136 20652 289142 20664
rect 579982 20652 579988 20664
rect 289136 20624 579988 20652
rect 289136 20612 289142 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 154390 20204 154396 20256
rect 154448 20244 154454 20256
rect 273254 20244 273260 20256
rect 154448 20216 273260 20244
rect 154448 20204 154454 20216
rect 273254 20204 273260 20216
rect 273312 20204 273318 20256
rect 153746 20136 153752 20188
rect 153804 20176 153810 20188
rect 280154 20176 280160 20188
rect 153804 20148 280160 20176
rect 153804 20136 153810 20148
rect 280154 20136 280160 20148
rect 280212 20136 280218 20188
rect 155770 20068 155776 20120
rect 155828 20108 155834 20120
rect 291194 20108 291200 20120
rect 155828 20080 291200 20108
rect 155828 20068 155834 20080
rect 291194 20068 291200 20080
rect 291252 20068 291258 20120
rect 161198 20000 161204 20052
rect 161256 20040 161262 20052
rect 372614 20040 372620 20052
rect 161256 20012 372620 20040
rect 161256 20000 161262 20012
rect 372614 20000 372620 20012
rect 372672 20000 372678 20052
rect 155678 19932 155684 19984
rect 155736 19972 155742 19984
rect 287054 19972 287060 19984
rect 155736 19944 287060 19972
rect 155736 19932 155742 19944
rect 287054 19932 287060 19944
rect 287112 19932 287118 19984
rect 287698 19932 287704 19984
rect 287756 19972 287762 19984
rect 518894 19972 518900 19984
rect 287756 19944 518900 19972
rect 287756 19932 287762 19944
rect 518894 19932 518900 19944
rect 518952 19932 518958 19984
rect 155862 18776 155868 18828
rect 155920 18816 155926 18828
rect 300854 18816 300860 18828
rect 155920 18788 300860 18816
rect 155920 18776 155926 18788
rect 300854 18776 300860 18788
rect 300912 18776 300918 18828
rect 176286 18708 176292 18760
rect 176344 18748 176350 18760
rect 522390 18748 522396 18760
rect 176344 18720 522396 18748
rect 176344 18708 176350 18720
rect 522390 18708 522396 18720
rect 522448 18708 522454 18760
rect 176378 18640 176384 18692
rect 176436 18680 176442 18692
rect 567194 18680 567200 18692
rect 176436 18652 567200 18680
rect 176436 18640 176442 18652
rect 567194 18640 567200 18652
rect 567252 18640 567258 18692
rect 177942 18572 177948 18624
rect 178000 18612 178006 18624
rect 574094 18612 574100 18624
rect 178000 18584 574100 18612
rect 178000 18572 178006 18584
rect 574094 18572 574100 18584
rect 574152 18572 574158 18624
rect 150618 17484 150624 17536
rect 150676 17524 150682 17536
rect 241514 17524 241520 17536
rect 150676 17496 241520 17524
rect 150676 17484 150682 17496
rect 241514 17484 241520 17496
rect 241572 17484 241578 17536
rect 165522 17416 165528 17468
rect 165580 17456 165586 17468
rect 418154 17456 418160 17468
rect 165580 17428 418160 17456
rect 165580 17416 165586 17428
rect 418154 17416 418160 17428
rect 418212 17416 418218 17468
rect 166810 17348 166816 17400
rect 166868 17388 166874 17400
rect 441614 17388 441620 17400
rect 166868 17360 441620 17388
rect 166868 17348 166874 17360
rect 441614 17348 441620 17360
rect 441672 17348 441678 17400
rect 168098 17280 168104 17332
rect 168156 17320 168162 17332
rect 445754 17320 445760 17332
rect 168156 17292 445760 17320
rect 168156 17280 168162 17292
rect 445754 17280 445760 17292
rect 445812 17280 445818 17332
rect 145558 17212 145564 17264
rect 145616 17252 145622 17264
rect 164878 17252 164884 17264
rect 145616 17224 164884 17252
rect 145616 17212 145622 17224
rect 164878 17212 164884 17224
rect 164936 17212 164942 17264
rect 169662 17212 169668 17264
rect 169720 17252 169726 17264
rect 477494 17252 477500 17264
rect 169720 17224 477500 17252
rect 169720 17212 169726 17224
rect 477494 17212 477500 17224
rect 477552 17212 477558 17264
rect 153010 16124 153016 16176
rect 153068 16164 153074 16176
rect 259546 16164 259552 16176
rect 153068 16136 259552 16164
rect 153068 16124 153074 16136
rect 259546 16124 259552 16136
rect 259604 16124 259610 16176
rect 161106 16056 161112 16108
rect 161164 16096 161170 16108
rect 361114 16096 361120 16108
rect 161164 16068 361120 16096
rect 161164 16056 161170 16068
rect 361114 16056 361120 16068
rect 361172 16056 361178 16108
rect 160094 15988 160100 16040
rect 160152 16028 160158 16040
rect 364610 16028 364616 16040
rect 160152 16000 364616 16028
rect 160152 15988 160158 16000
rect 364610 15988 364616 16000
rect 364668 15988 364674 16040
rect 164142 15920 164148 15972
rect 164200 15960 164206 15972
rect 397730 15960 397736 15972
rect 164200 15932 397736 15960
rect 164200 15920 164206 15932
rect 397730 15920 397736 15932
rect 397788 15920 397794 15972
rect 400858 15920 400864 15972
rect 400916 15960 400922 15972
rect 478874 15960 478880 15972
rect 400916 15932 478880 15960
rect 400916 15920 400922 15932
rect 478874 15920 478880 15932
rect 478932 15920 478938 15972
rect 165338 15852 165344 15904
rect 165396 15892 165402 15904
rect 420914 15892 420920 15904
rect 165396 15864 420920 15892
rect 165396 15852 165402 15864
rect 420914 15852 420920 15864
rect 420972 15852 420978 15904
rect 153930 14696 153936 14748
rect 153988 14736 153994 14748
rect 272426 14736 272432 14748
rect 153988 14708 272432 14736
rect 153988 14696 153994 14708
rect 272426 14696 272432 14708
rect 272484 14696 272490 14748
rect 156782 14628 156788 14680
rect 156840 14668 156846 14680
rect 314654 14668 314660 14680
rect 156840 14640 314660 14668
rect 156840 14628 156846 14640
rect 314654 14628 314660 14640
rect 314712 14628 314718 14680
rect 179322 14560 179328 14612
rect 179380 14600 179386 14612
rect 394234 14600 394240 14612
rect 179380 14572 394240 14600
rect 179380 14560 179386 14572
rect 394234 14560 394240 14572
rect 394292 14560 394298 14612
rect 164050 14492 164056 14544
rect 164108 14532 164114 14544
rect 407206 14532 407212 14544
rect 164108 14504 407212 14532
rect 164108 14492 164114 14504
rect 407206 14492 407212 14504
rect 407264 14492 407270 14544
rect 171870 14424 171876 14476
rect 171928 14464 171934 14476
rect 503714 14464 503720 14476
rect 171928 14436 503720 14464
rect 171928 14424 171934 14436
rect 503714 14424 503720 14436
rect 503772 14424 503778 14476
rect 153838 13336 153844 13388
rect 153896 13376 153902 13388
rect 276014 13376 276020 13388
rect 153896 13348 276020 13376
rect 153896 13336 153902 13348
rect 276014 13336 276020 13348
rect 276072 13336 276078 13388
rect 158530 13268 158536 13320
rect 158588 13308 158594 13320
rect 324406 13308 324412 13320
rect 158588 13280 324412 13308
rect 158588 13268 158594 13280
rect 324406 13268 324412 13280
rect 324464 13268 324470 13320
rect 178770 13200 178776 13252
rect 178828 13240 178834 13252
rect 400858 13240 400864 13252
rect 178828 13212 400864 13240
rect 178828 13200 178834 13212
rect 400858 13200 400864 13212
rect 400916 13200 400922 13252
rect 165430 13132 165436 13184
rect 165488 13172 165494 13184
rect 414290 13172 414296 13184
rect 165488 13144 414296 13172
rect 165488 13132 165494 13144
rect 414290 13132 414296 13144
rect 414348 13132 414354 13184
rect 172054 13064 172060 13116
rect 172112 13104 172118 13116
rect 511258 13104 511264 13116
rect 172112 13076 511264 13104
rect 172112 13064 172118 13076
rect 511258 13064 511264 13076
rect 511316 13064 511322 13116
rect 150894 11908 150900 11960
rect 150952 11948 150958 11960
rect 245194 11948 245200 11960
rect 150952 11920 245200 11948
rect 150952 11908 150958 11920
rect 245194 11908 245200 11920
rect 245252 11908 245258 11960
rect 162670 11840 162676 11892
rect 162728 11880 162734 11892
rect 386690 11880 386696 11892
rect 162728 11852 386696 11880
rect 162728 11840 162734 11852
rect 386690 11840 386696 11852
rect 386748 11840 386754 11892
rect 165614 11772 165620 11824
rect 165672 11812 165678 11824
rect 439130 11812 439136 11824
rect 165672 11784 439136 11812
rect 165672 11772 165678 11784
rect 439130 11772 439136 11784
rect 439188 11772 439194 11824
rect 175090 11704 175096 11756
rect 175148 11744 175154 11756
rect 548610 11744 548616 11756
rect 175148 11716 548616 11744
rect 175148 11704 175154 11716
rect 548610 11704 548616 11716
rect 548668 11704 548674 11756
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 152458 10548 152464 10600
rect 152516 10588 152522 10600
rect 258258 10588 258264 10600
rect 152516 10560 258264 10588
rect 152516 10548 152522 10560
rect 258258 10548 258264 10560
rect 258316 10548 258322 10600
rect 156690 10480 156696 10532
rect 156748 10520 156754 10532
rect 307938 10520 307944 10532
rect 156748 10492 307944 10520
rect 156748 10480 156754 10492
rect 307938 10480 307944 10492
rect 307996 10480 308002 10532
rect 162486 10412 162492 10464
rect 162544 10452 162550 10464
rect 385954 10452 385960 10464
rect 162544 10424 385960 10452
rect 162544 10412 162550 10424
rect 385954 10412 385960 10424
rect 386012 10412 386018 10464
rect 162762 10344 162768 10396
rect 162820 10384 162826 10396
rect 390646 10384 390652 10396
rect 162820 10356 390652 10384
rect 162820 10344 162826 10356
rect 390646 10344 390652 10356
rect 390704 10344 390710 10396
rect 87506 10276 87512 10328
rect 87564 10316 87570 10328
rect 138106 10316 138112 10328
rect 87564 10288 138112 10316
rect 87564 10276 87570 10288
rect 138106 10276 138112 10288
rect 138164 10276 138170 10328
rect 170950 10276 170956 10328
rect 171008 10316 171014 10328
rect 493042 10316 493048 10328
rect 171008 10288 493048 10316
rect 171008 10276 171014 10288
rect 493042 10276 493048 10288
rect 493100 10276 493106 10328
rect 151170 9256 151176 9308
rect 151228 9296 151234 9308
rect 234706 9296 234712 9308
rect 151228 9268 234712 9296
rect 151228 9256 151234 9268
rect 234706 9256 234712 9268
rect 234764 9256 234770 9308
rect 158622 9188 158628 9240
rect 158680 9228 158686 9240
rect 329190 9228 329196 9240
rect 158680 9200 329196 9228
rect 158680 9188 158686 9200
rect 329190 9188 329196 9200
rect 329248 9188 329254 9240
rect 161382 9120 161388 9172
rect 161440 9160 161446 9172
rect 365806 9160 365812 9172
rect 161440 9132 365812 9160
rect 161440 9120 161446 9132
rect 365806 9120 365812 9132
rect 365864 9120 365870 9172
rect 166902 9052 166908 9104
rect 166960 9092 166966 9104
rect 432046 9092 432052 9104
rect 166960 9064 432052 9092
rect 166960 9052 166966 9064
rect 432046 9052 432052 9064
rect 432104 9052 432110 9104
rect 176470 8984 176476 9036
rect 176528 9024 176534 9036
rect 556154 9024 556160 9036
rect 176528 8996 556160 9024
rect 176528 8984 176534 8996
rect 556154 8984 556160 8996
rect 556212 8984 556218 9036
rect 105722 8916 105728 8968
rect 105780 8956 105786 8968
rect 139854 8956 139860 8968
rect 105780 8928 139860 8956
rect 105780 8916 105786 8928
rect 139854 8916 139860 8928
rect 139912 8916 139918 8968
rect 143534 8916 143540 8968
rect 143592 8956 143598 8968
rect 151906 8956 151912 8968
rect 143592 8928 151912 8956
rect 143592 8916 143598 8928
rect 151906 8916 151912 8928
rect 151964 8916 151970 8968
rect 185578 8916 185584 8968
rect 185636 8956 185642 8968
rect 580994 8956 581000 8968
rect 185636 8928 581000 8956
rect 185636 8916 185642 8928
rect 580994 8916 581000 8928
rect 581052 8916 581058 8968
rect 149146 7760 149152 7812
rect 149204 7800 149210 7812
rect 227530 7800 227536 7812
rect 149204 7772 227536 7800
rect 149204 7760 149210 7772
rect 227530 7760 227536 7772
rect 227588 7760 227594 7812
rect 160002 7692 160008 7744
rect 160060 7732 160066 7744
rect 350442 7732 350448 7744
rect 160060 7704 350448 7732
rect 160060 7692 160066 7704
rect 350442 7692 350448 7704
rect 350500 7692 350506 7744
rect 168282 7624 168288 7676
rect 168340 7664 168346 7676
rect 453390 7664 453396 7676
rect 168340 7636 453396 7664
rect 168340 7624 168346 7636
rect 453390 7624 453396 7636
rect 453448 7624 453454 7676
rect 30098 7556 30104 7608
rect 30156 7596 30162 7608
rect 134150 7596 134156 7608
rect 30156 7568 134156 7596
rect 30156 7556 30162 7568
rect 134150 7556 134156 7568
rect 134208 7556 134214 7608
rect 175182 7556 175188 7608
rect 175240 7596 175246 7608
rect 545482 7596 545488 7608
rect 175240 7568 545488 7596
rect 175240 7556 175246 7568
rect 545482 7556 545488 7568
rect 545540 7556 545546 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 17218 6848 17224 6860
rect 3476 6820 17224 6848
rect 3476 6808 3482 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 576118 6808 576124 6860
rect 576176 6848 576182 6860
rect 580166 6848 580172 6860
rect 576176 6820 580172 6848
rect 576176 6808 576182 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 156414 6400 156420 6452
rect 156472 6440 156478 6452
rect 316218 6440 316224 6452
rect 156472 6412 316224 6440
rect 156472 6400 156478 6412
rect 316218 6400 316224 6412
rect 316276 6400 316282 6452
rect 161290 6332 161296 6384
rect 161348 6372 161354 6384
rect 371694 6372 371700 6384
rect 161348 6344 371700 6372
rect 161348 6332 161354 6344
rect 371694 6332 371700 6344
rect 371752 6332 371758 6384
rect 169754 6264 169760 6316
rect 169812 6304 169818 6316
rect 482830 6304 482836 6316
rect 169812 6276 482836 6304
rect 169812 6264 169818 6276
rect 482830 6264 482836 6276
rect 482888 6264 482894 6316
rect 176562 6196 176568 6248
rect 176620 6236 176626 6248
rect 558546 6236 558552 6248
rect 176620 6208 558552 6236
rect 176620 6196 176626 6208
rect 558546 6196 558552 6208
rect 558604 6196 558610 6248
rect 175826 6128 175832 6180
rect 175884 6168 175890 6180
rect 563238 6168 563244 6180
rect 175884 6140 563244 6168
rect 175884 6128 175890 6140
rect 563238 6128 563244 6140
rect 563296 6128 563302 6180
rect 152090 4972 152096 5024
rect 152148 5012 152154 5024
rect 266538 5012 266544 5024
rect 152148 4984 266544 5012
rect 152148 4972 152154 4984
rect 266538 4972 266544 4984
rect 266596 4972 266602 5024
rect 162578 4904 162584 4956
rect 162636 4944 162642 4956
rect 378870 4944 378876 4956
rect 162636 4916 378876 4944
rect 162636 4904 162642 4916
rect 378870 4904 378876 4916
rect 378928 4904 378934 4956
rect 170398 4836 170404 4888
rect 170456 4876 170462 4888
rect 486326 4876 486332 4888
rect 170456 4848 486332 4876
rect 170456 4836 170462 4848
rect 486326 4836 486332 4848
rect 486384 4836 486390 4888
rect 173894 4768 173900 4820
rect 173952 4808 173958 4820
rect 541986 4808 541992 4820
rect 173952 4780 541992 4808
rect 173952 4768 173958 4780
rect 541986 4768 541992 4780
rect 542044 4768 542050 4820
rect 142798 4156 142804 4208
rect 142856 4196 142862 4208
rect 143534 4196 143540 4208
rect 142856 4168 143540 4196
rect 142856 4156 142862 4168
rect 143534 4156 143540 4168
rect 143592 4156 143598 4208
rect 566 4088 572 4140
rect 624 4128 630 4140
rect 7558 4128 7564 4140
rect 624 4100 7564 4128
rect 624 4088 630 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 17310 4128 17316 4140
rect 15988 4100 17316 4128
rect 15988 4088 15994 4100
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 73798 4088 73804 4140
rect 73856 4128 73862 4140
rect 75178 4128 75184 4140
rect 73856 4100 75184 4128
rect 73856 4088 73862 4100
rect 75178 4088 75184 4100
rect 75236 4088 75242 4140
rect 127618 4088 127624 4140
rect 127676 4128 127682 4140
rect 134518 4128 134524 4140
rect 127676 4100 134524 4128
rect 127676 4088 127682 4100
rect 134518 4088 134524 4100
rect 134576 4088 134582 4140
rect 146938 4088 146944 4140
rect 146996 4128 147002 4140
rect 147398 4128 147404 4140
rect 146996 4100 147404 4128
rect 146996 4088 147002 4100
rect 147398 4088 147404 4100
rect 147456 4088 147462 4140
rect 169018 4088 169024 4140
rect 169076 4128 169082 4140
rect 173158 4128 173164 4140
rect 169076 4100 173164 4128
rect 169076 4088 169082 4100
rect 173158 4088 173164 4100
rect 173216 4088 173222 4140
rect 196618 4088 196624 4140
rect 196676 4128 196682 4140
rect 200298 4128 200304 4140
rect 196676 4100 200304 4128
rect 196676 4088 196682 4100
rect 200298 4088 200304 4100
rect 200356 4088 200362 4140
rect 301590 4088 301596 4140
rect 301648 4128 301654 4140
rect 309042 4128 309048 4140
rect 301648 4100 309048 4128
rect 301648 4088 301654 4100
rect 309042 4088 309048 4100
rect 309100 4088 309106 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 317322 4128 317328 4140
rect 315356 4100 317328 4128
rect 315356 4088 315362 4100
rect 317322 4088 317328 4100
rect 317380 4088 317386 4140
rect 324958 4088 324964 4140
rect 325016 4128 325022 4140
rect 326798 4128 326804 4140
rect 325016 4100 326804 4128
rect 325016 4088 325022 4100
rect 326798 4088 326804 4100
rect 326856 4088 326862 4140
rect 382918 4088 382924 4140
rect 382976 4128 382982 4140
rect 384758 4128 384764 4140
rect 382976 4100 384764 4128
rect 382976 4088 382982 4100
rect 384758 4088 384764 4100
rect 384816 4088 384822 4140
rect 450538 4088 450544 4140
rect 450596 4128 450602 4140
rect 452102 4128 452108 4140
rect 450596 4100 452108 4128
rect 450596 4088 450602 4100
rect 452102 4088 452108 4100
rect 452160 4088 452166 4140
rect 489178 4088 489184 4140
rect 489236 4128 489242 4140
rect 491110 4128 491116 4140
rect 489236 4100 491116 4128
rect 489236 4088 489242 4100
rect 491110 4088 491116 4100
rect 491168 4088 491174 4140
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 8938 4060 8944 4072
rect 1728 4032 8944 4060
rect 1728 4020 1734 4032
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 147306 4020 147312 4072
rect 147364 4060 147370 4072
rect 150710 4060 150716 4072
rect 147364 4032 150716 4060
rect 147364 4020 147370 4032
rect 150710 4020 150716 4032
rect 150768 4020 150774 4072
rect 151814 4020 151820 4072
rect 151872 4060 151878 4072
rect 153010 4060 153016 4072
rect 151872 4032 153016 4060
rect 151872 4020 151878 4032
rect 153010 4020 153016 4032
rect 153068 4020 153074 4072
rect 130838 3952 130844 4004
rect 130896 3992 130902 4004
rect 144730 3992 144736 4004
rect 130896 3964 144736 3992
rect 130896 3952 130902 3964
rect 144730 3952 144736 3964
rect 144788 3952 144794 4004
rect 149698 3952 149704 4004
rect 149756 3992 149762 4004
rect 157794 3992 157800 4004
rect 149756 3964 157800 3992
rect 149756 3952 149762 3964
rect 157794 3952 157800 3964
rect 157852 3952 157858 4004
rect 45922 3884 45928 3936
rect 45980 3924 45986 3936
rect 46198 3924 46204 3936
rect 45980 3896 46204 3924
rect 45980 3884 45986 3896
rect 46198 3884 46204 3896
rect 46256 3884 46262 3936
rect 124674 3884 124680 3936
rect 124732 3924 124738 3936
rect 140866 3924 140872 3936
rect 124732 3896 140872 3924
rect 124732 3884 124738 3896
rect 140866 3884 140872 3896
rect 140924 3884 140930 3936
rect 149790 3884 149796 3936
rect 149848 3924 149854 3936
rect 156598 3924 156604 3936
rect 149848 3896 156604 3924
rect 149848 3884 149854 3896
rect 156598 3884 156604 3896
rect 156656 3884 156662 3936
rect 156690 3884 156696 3936
rect 156748 3924 156754 3936
rect 170766 3924 170772 3936
rect 156748 3896 170772 3924
rect 156748 3884 156754 3896
rect 170766 3884 170772 3896
rect 170824 3884 170830 3936
rect 112806 3816 112812 3868
rect 112864 3856 112870 3868
rect 117406 3856 117412 3868
rect 112864 3828 117412 3856
rect 112864 3816 112870 3828
rect 117406 3816 117412 3828
rect 117464 3816 117470 3868
rect 125870 3816 125876 3868
rect 125928 3856 125934 3868
rect 129918 3856 129924 3868
rect 125928 3828 129924 3856
rect 125928 3816 125934 3828
rect 129918 3816 129924 3828
rect 129976 3816 129982 3868
rect 130746 3816 130752 3868
rect 130804 3856 130810 3868
rect 162486 3856 162492 3868
rect 130804 3828 162492 3856
rect 130804 3816 130810 3828
rect 162486 3816 162492 3828
rect 162544 3816 162550 3868
rect 91554 3748 91560 3800
rect 91612 3788 91618 3800
rect 139486 3788 139492 3800
rect 91612 3760 139492 3788
rect 91612 3748 91618 3760
rect 139486 3748 139492 3760
rect 139544 3748 139550 3800
rect 147214 3748 147220 3800
rect 147272 3788 147278 3800
rect 163682 3788 163688 3800
rect 147272 3760 163688 3788
rect 147272 3748 147278 3760
rect 163682 3748 163688 3760
rect 163740 3748 163746 3800
rect 164712 3760 171134 3788
rect 85666 3680 85672 3732
rect 85724 3720 85730 3732
rect 127618 3720 127624 3732
rect 85724 3692 127624 3720
rect 85724 3680 85730 3692
rect 127618 3680 127624 3692
rect 127676 3680 127682 3732
rect 129826 3720 129832 3732
rect 127820 3692 129832 3720
rect 66714 3612 66720 3664
rect 66772 3652 66778 3664
rect 72418 3652 72424 3664
rect 66772 3624 72424 3652
rect 66772 3612 66778 3624
rect 72418 3612 72424 3624
rect 72476 3612 72482 3664
rect 83274 3612 83280 3664
rect 83332 3652 83338 3664
rect 127710 3652 127716 3664
rect 83332 3624 127716 3652
rect 83332 3612 83338 3624
rect 127710 3612 127716 3624
rect 127768 3612 127774 3664
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 21358 3584 21364 3596
rect 19484 3556 21364 3584
rect 19484 3544 19490 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 44174 3544 44180 3596
rect 44232 3584 44238 3596
rect 45094 3584 45100 3596
rect 44232 3556 45100 3584
rect 44232 3544 44238 3556
rect 45094 3544 45100 3556
rect 45152 3544 45158 3596
rect 51350 3544 51356 3596
rect 51408 3584 51414 3596
rect 54478 3584 54484 3596
rect 51408 3556 54484 3584
rect 51408 3544 51414 3556
rect 54478 3544 54484 3556
rect 54536 3544 54542 3596
rect 59630 3544 59636 3596
rect 59688 3584 59694 3596
rect 64138 3584 64144 3596
rect 59688 3556 64144 3584
rect 59688 3544 59694 3556
rect 64138 3544 64144 3556
rect 64196 3544 64202 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 127820 3584 127848 3692
rect 129826 3680 129832 3692
rect 129884 3680 129890 3732
rect 138198 3720 138204 3732
rect 132466 3692 138204 3720
rect 127894 3612 127900 3664
rect 127952 3652 127958 3664
rect 132466 3652 132494 3692
rect 138198 3680 138204 3692
rect 138256 3680 138262 3732
rect 147122 3680 147128 3732
rect 147180 3720 147186 3732
rect 150618 3720 150624 3732
rect 147180 3692 150624 3720
rect 147180 3680 147186 3692
rect 150618 3680 150624 3692
rect 150676 3680 150682 3732
rect 150710 3680 150716 3732
rect 150768 3720 150774 3732
rect 164510 3720 164516 3732
rect 150768 3692 164516 3720
rect 150768 3680 150774 3692
rect 164510 3680 164516 3692
rect 164568 3680 164574 3732
rect 127952 3624 132494 3652
rect 127952 3612 127958 3624
rect 137646 3612 137652 3664
rect 137704 3652 137710 3664
rect 138658 3652 138664 3664
rect 137704 3624 138664 3652
rect 137704 3612 137710 3624
rect 138658 3612 138664 3624
rect 138716 3612 138722 3664
rect 147030 3612 147036 3664
rect 147088 3652 147094 3664
rect 149514 3652 149520 3664
rect 147088 3624 149520 3652
rect 147088 3612 147094 3624
rect 149514 3612 149520 3624
rect 149572 3612 149578 3664
rect 151078 3612 151084 3664
rect 151136 3652 151142 3664
rect 164712 3652 164740 3760
rect 166074 3720 166080 3732
rect 151136 3624 164740 3652
rect 164804 3692 166080 3720
rect 151136 3612 151142 3624
rect 69164 3556 127848 3584
rect 69164 3544 69170 3556
rect 128170 3544 128176 3596
rect 128228 3584 128234 3596
rect 130378 3584 130384 3596
rect 128228 3556 130384 3584
rect 128228 3544 128234 3556
rect 130378 3544 130384 3556
rect 130436 3544 130442 3596
rect 130930 3544 130936 3596
rect 130988 3584 130994 3596
rect 164804 3584 164832 3692
rect 166074 3680 166080 3692
rect 166132 3680 166138 3732
rect 171106 3652 171134 3760
rect 184198 3748 184204 3800
rect 184256 3788 184262 3800
rect 210970 3788 210976 3800
rect 184256 3760 210976 3788
rect 184256 3748 184262 3760
rect 210970 3748 210976 3760
rect 211028 3748 211034 3800
rect 211798 3748 211804 3800
rect 211856 3788 211862 3800
rect 211856 3760 219434 3788
rect 211856 3748 211862 3760
rect 181438 3680 181444 3732
rect 181496 3720 181502 3732
rect 212166 3720 212172 3732
rect 181496 3692 212172 3720
rect 181496 3680 181502 3692
rect 212166 3680 212172 3692
rect 212224 3680 212230 3732
rect 219406 3720 219434 3760
rect 234614 3748 234620 3800
rect 234672 3788 234678 3800
rect 235810 3788 235816 3800
rect 234672 3760 235816 3788
rect 234672 3748 234678 3760
rect 235810 3748 235816 3760
rect 235868 3748 235874 3800
rect 247586 3720 247592 3732
rect 219406 3692 247592 3720
rect 247586 3680 247592 3692
rect 247644 3680 247650 3732
rect 423766 3680 423772 3732
rect 423824 3720 423830 3732
rect 424962 3720 424968 3732
rect 423824 3692 424968 3720
rect 423824 3680 423830 3692
rect 424962 3680 424968 3692
rect 425020 3680 425026 3732
rect 171962 3652 171968 3664
rect 171106 3624 171968 3652
rect 171962 3612 171968 3624
rect 172020 3612 172026 3664
rect 189810 3612 189816 3664
rect 189868 3652 189874 3664
rect 193214 3652 193220 3664
rect 189868 3624 193220 3652
rect 189868 3612 189874 3624
rect 193214 3612 193220 3624
rect 193272 3612 193278 3664
rect 203702 3612 203708 3664
rect 203760 3652 203766 3664
rect 240502 3652 240508 3664
rect 203760 3624 240508 3652
rect 203760 3612 203766 3624
rect 240502 3612 240508 3624
rect 240560 3612 240566 3664
rect 247678 3612 247684 3664
rect 247736 3652 247742 3664
rect 254670 3652 254676 3664
rect 247736 3624 254676 3652
rect 247736 3612 247742 3624
rect 254670 3612 254676 3624
rect 254728 3612 254734 3664
rect 261478 3612 261484 3664
rect 261536 3652 261542 3664
rect 262950 3652 262956 3664
rect 261536 3624 262956 3652
rect 261536 3612 261542 3624
rect 262950 3612 262956 3624
rect 263008 3612 263014 3664
rect 299566 3612 299572 3664
rect 299624 3652 299630 3664
rect 300762 3652 300768 3664
rect 299624 3624 300768 3652
rect 299624 3612 299630 3624
rect 300762 3612 300768 3624
rect 300820 3612 300826 3664
rect 311158 3612 311164 3664
rect 311216 3652 311222 3664
rect 312630 3652 312636 3664
rect 311216 3624 312636 3652
rect 311216 3612 311222 3624
rect 312630 3612 312636 3624
rect 312688 3612 312694 3664
rect 130988 3556 164832 3584
rect 130988 3544 130994 3556
rect 164878 3544 164884 3596
rect 164936 3584 164942 3596
rect 168374 3584 168380 3596
rect 164936 3556 168380 3584
rect 164936 3544 164942 3556
rect 168374 3544 168380 3556
rect 168432 3544 168438 3596
rect 173250 3544 173256 3596
rect 173308 3584 173314 3596
rect 177850 3584 177856 3596
rect 173308 3556 177856 3584
rect 173308 3544 173314 3556
rect 177850 3544 177856 3556
rect 177908 3544 177914 3596
rect 180058 3544 180064 3596
rect 180116 3544 180122 3596
rect 181530 3544 181536 3596
rect 181588 3584 181594 3596
rect 182542 3584 182548 3596
rect 181588 3556 182548 3584
rect 181588 3544 181594 3556
rect 182542 3544 182548 3556
rect 182600 3544 182606 3596
rect 183002 3544 183008 3596
rect 183060 3584 183066 3596
rect 190822 3584 190828 3596
rect 183060 3556 190828 3584
rect 183060 3544 183066 3556
rect 190822 3544 190828 3556
rect 190880 3544 190886 3596
rect 193858 3544 193864 3596
rect 193916 3584 193922 3596
rect 196802 3584 196808 3596
rect 193916 3556 196808 3584
rect 193916 3544 193922 3556
rect 196802 3544 196808 3556
rect 196860 3544 196866 3596
rect 206278 3544 206284 3596
rect 206336 3584 206342 3596
rect 403618 3584 403624 3596
rect 206336 3556 403624 3584
rect 206336 3544 206342 3556
rect 403618 3544 403624 3556
rect 403676 3544 403682 3596
rect 407114 3544 407120 3596
rect 407172 3584 407178 3596
rect 408402 3584 408408 3596
rect 407172 3556 408408 3584
rect 407172 3544 407178 3556
rect 408402 3544 408408 3556
rect 408460 3544 408466 3596
rect 410518 3544 410524 3596
rect 410576 3584 410582 3596
rect 411898 3584 411904 3596
rect 410576 3556 411904 3584
rect 410576 3544 410582 3556
rect 411898 3544 411904 3556
rect 411956 3544 411962 3596
rect 418798 3544 418804 3596
rect 418856 3584 418862 3596
rect 420178 3584 420184 3596
rect 418856 3556 420184 3584
rect 418856 3544 418862 3556
rect 420178 3544 420184 3556
rect 420236 3544 420242 3596
rect 422938 3544 422944 3596
rect 422996 3584 423002 3596
rect 423766 3584 423772 3596
rect 422996 3556 423772 3584
rect 422996 3544 423002 3556
rect 423766 3544 423772 3556
rect 423824 3544 423830 3596
rect 431954 3544 431960 3596
rect 432012 3584 432018 3596
rect 433242 3584 433248 3596
rect 432012 3556 433248 3584
rect 432012 3544 432018 3556
rect 433242 3544 433248 3556
rect 433300 3544 433306 3596
rect 440234 3544 440240 3596
rect 440292 3584 440298 3596
rect 441522 3584 441528 3596
rect 440292 3556 441528 3584
rect 440292 3544 440298 3556
rect 441522 3544 441528 3556
rect 441580 3544 441586 3596
rect 446398 3544 446404 3596
rect 446456 3584 446462 3596
rect 447410 3584 447416 3596
rect 446456 3556 447416 3584
rect 446456 3544 446462 3556
rect 447410 3544 447416 3556
rect 447468 3544 447474 3596
rect 448606 3544 448612 3596
rect 448664 3584 448670 3596
rect 449802 3584 449808 3596
rect 448664 3556 449808 3584
rect 448664 3544 448670 3556
rect 449802 3544 449808 3556
rect 449860 3544 449866 3596
rect 453298 3544 453304 3596
rect 453356 3584 453362 3596
rect 497090 3584 497096 3596
rect 453356 3556 497096 3584
rect 453356 3544 453362 3556
rect 497090 3544 497096 3556
rect 497148 3544 497154 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 576302 3584 576308 3596
rect 574796 3556 576308 3584
rect 574796 3544 574802 3556
rect 576302 3544 576308 3556
rect 576360 3544 576366 3596
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6512 3488 123340 3516
rect 6512 3476 6518 3488
rect 8754 3408 8760 3460
rect 8812 3448 8818 3460
rect 10318 3448 10324 3460
rect 8812 3420 10324 3448
rect 8812 3408 8818 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 18598 3448 18604 3460
rect 17092 3420 18604 3448
rect 17092 3408 17098 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 27614 3408 27620 3460
rect 27672 3448 27678 3460
rect 28534 3448 28540 3460
rect 27672 3420 28540 3448
rect 27672 3408 27678 3420
rect 28534 3408 28540 3420
rect 28592 3408 28598 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 45922 3448 45928 3460
rect 33652 3420 45928 3448
rect 33652 3408 33658 3420
rect 45922 3408 45928 3420
rect 45980 3408 45986 3460
rect 52454 3408 52460 3460
rect 52512 3448 52518 3460
rect 53374 3448 53380 3460
rect 52512 3420 53380 3448
rect 52512 3408 52518 3420
rect 53374 3408 53380 3420
rect 53432 3408 53438 3460
rect 56042 3408 56048 3460
rect 56100 3448 56106 3460
rect 57238 3448 57244 3460
rect 56100 3420 57244 3448
rect 56100 3408 56106 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 60734 3408 60740 3460
rect 60792 3448 60798 3460
rect 61654 3448 61660 3460
rect 60792 3420 61660 3448
rect 60792 3408 60798 3420
rect 61654 3408 61660 3420
rect 61712 3408 61718 3460
rect 65518 3408 65524 3460
rect 65576 3448 65582 3460
rect 65576 3420 122834 3448
rect 65576 3408 65582 3420
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 122806 3312 122834 3420
rect 123312 3380 123340 3488
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124950 3516 124956 3528
rect 123536 3488 124956 3516
rect 123536 3476 123542 3488
rect 124950 3476 124956 3488
rect 125008 3476 125014 3528
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128446 3516 128452 3528
rect 127032 3488 128452 3516
rect 127032 3476 127038 3488
rect 128446 3476 128452 3488
rect 128504 3476 128510 3528
rect 175458 3516 175464 3528
rect 150820 3488 175464 3516
rect 137278 3448 137284 3460
rect 132466 3420 137284 3448
rect 131758 3380 131764 3392
rect 123312 3352 131764 3380
rect 131758 3340 131764 3352
rect 131816 3340 131822 3392
rect 132466 3312 132494 3420
rect 137278 3408 137284 3420
rect 137336 3408 137342 3460
rect 148318 3408 148324 3460
rect 148376 3448 148382 3460
rect 150820 3448 150848 3488
rect 175458 3476 175464 3488
rect 175516 3476 175522 3528
rect 180076 3516 180104 3544
rect 458082 3516 458088 3528
rect 180076 3488 458088 3516
rect 458082 3476 458088 3488
rect 458140 3476 458146 3528
rect 468478 3476 468484 3528
rect 468536 3516 468542 3528
rect 469858 3516 469864 3528
rect 468536 3488 469864 3516
rect 468536 3476 468542 3488
rect 469858 3476 469864 3488
rect 469916 3476 469922 3528
rect 472618 3476 472624 3528
rect 472676 3516 472682 3528
rect 473446 3516 473452 3528
rect 472676 3488 473452 3516
rect 472676 3476 472682 3488
rect 473446 3476 473452 3488
rect 473504 3476 473510 3528
rect 486418 3476 486424 3528
rect 486476 3516 486482 3528
rect 487614 3516 487620 3528
rect 486476 3488 487620 3516
rect 486476 3476 486482 3488
rect 487614 3476 487620 3488
rect 487672 3476 487678 3528
rect 504358 3476 504364 3528
rect 504416 3516 504422 3528
rect 505370 3516 505376 3528
rect 504416 3488 505376 3516
rect 504416 3476 504422 3488
rect 505370 3476 505376 3488
rect 505428 3476 505434 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 509878 3476 509884 3528
rect 509936 3516 509942 3528
rect 518342 3516 518348 3528
rect 509936 3488 518348 3516
rect 509936 3476 509942 3488
rect 518342 3476 518348 3488
rect 518400 3476 518406 3528
rect 527910 3476 527916 3528
rect 527968 3516 527974 3528
rect 533706 3516 533712 3528
rect 527968 3488 533712 3516
rect 527968 3476 527974 3488
rect 533706 3476 533712 3488
rect 533764 3476 533770 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 545758 3476 545764 3528
rect 545816 3516 545822 3528
rect 551462 3516 551468 3528
rect 545816 3488 551468 3516
rect 545816 3476 545822 3488
rect 551462 3476 551468 3488
rect 551520 3476 551526 3528
rect 558178 3476 558184 3528
rect 558236 3516 558242 3528
rect 559742 3516 559748 3528
rect 558236 3488 559748 3516
rect 558236 3476 558242 3488
rect 559742 3476 559748 3488
rect 559800 3476 559806 3528
rect 563698 3476 563704 3528
rect 563756 3516 563762 3528
rect 565630 3516 565636 3528
rect 563756 3488 565636 3516
rect 563756 3476 563762 3488
rect 565630 3476 565636 3488
rect 565688 3476 565694 3528
rect 567838 3476 567844 3528
rect 567896 3516 567902 3528
rect 569126 3516 569132 3528
rect 567896 3488 569132 3516
rect 567896 3476 567902 3488
rect 569126 3476 569132 3488
rect 569184 3476 569190 3528
rect 571978 3476 571984 3528
rect 572036 3516 572042 3528
rect 573910 3516 573916 3528
rect 572036 3488 573916 3516
rect 572036 3476 572042 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 176654 3448 176660 3460
rect 148376 3420 150848 3448
rect 151786 3420 176660 3448
rect 148376 3408 148382 3420
rect 147398 3340 147404 3392
rect 147456 3380 147462 3392
rect 151786 3380 151814 3420
rect 176654 3408 176660 3420
rect 176712 3408 176718 3460
rect 178678 3408 178684 3460
rect 178736 3448 178742 3460
rect 468662 3448 468668 3460
rect 178736 3420 468668 3448
rect 178736 3408 178742 3420
rect 468662 3408 468668 3420
rect 468720 3408 468726 3460
rect 480898 3408 480904 3460
rect 480956 3448 480962 3460
rect 521838 3448 521844 3460
rect 480956 3420 521844 3448
rect 480956 3408 480962 3420
rect 521838 3408 521844 3420
rect 521896 3408 521902 3460
rect 522390 3408 522396 3460
rect 522448 3448 522454 3460
rect 560846 3448 560852 3460
rect 522448 3420 560852 3448
rect 522448 3408 522454 3420
rect 560846 3408 560852 3420
rect 560904 3408 560910 3460
rect 560938 3408 560944 3460
rect 560996 3448 561002 3460
rect 572714 3448 572720 3460
rect 560996 3420 572720 3448
rect 560996 3408 561002 3420
rect 572714 3408 572720 3420
rect 572772 3408 572778 3460
rect 147456 3352 151814 3380
rect 147456 3340 147462 3352
rect 275278 3340 275284 3392
rect 275336 3380 275342 3392
rect 277118 3380 277124 3392
rect 275336 3352 277124 3380
rect 275336 3340 275342 3352
rect 277118 3340 277124 3352
rect 277176 3340 277182 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 340874 3340 340880 3392
rect 340932 3380 340938 3392
rect 342162 3380 342168 3392
rect 340932 3352 342168 3380
rect 340932 3340 340938 3352
rect 342162 3340 342168 3352
rect 342220 3340 342226 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 364978 3340 364984 3392
rect 365036 3380 365042 3392
rect 367002 3380 367008 3392
rect 365036 3352 367008 3380
rect 365036 3340 365042 3352
rect 367002 3340 367008 3352
rect 367060 3340 367066 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 414658 3340 414664 3392
rect 414716 3380 414722 3392
rect 416682 3380 416688 3392
rect 414716 3352 416688 3380
rect 414716 3340 414722 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 122806 3284 132494 3312
rect 38378 3136 38384 3188
rect 38436 3176 38442 3188
rect 39298 3176 39304 3188
rect 38436 3148 39304 3176
rect 38436 3136 38442 3148
rect 39298 3136 39304 3148
rect 39356 3136 39362 3188
rect 148410 3136 148416 3188
rect 148468 3176 148474 3188
rect 154206 3176 154212 3188
rect 148468 3148 154212 3176
rect 148468 3136 148474 3148
rect 154206 3136 154212 3148
rect 154264 3136 154270 3188
rect 171778 3136 171784 3188
rect 171836 3176 171842 3188
rect 174262 3176 174268 3188
rect 171836 3148 174268 3176
rect 171836 3136 171842 3148
rect 174262 3136 174268 3148
rect 174320 3136 174326 3188
rect 200758 3136 200764 3188
rect 200816 3176 200822 3188
rect 203886 3176 203892 3188
rect 200816 3148 203892 3176
rect 200816 3136 200822 3148
rect 203886 3136 203892 3148
rect 203944 3136 203950 3188
rect 297358 3136 297364 3188
rect 297416 3176 297422 3188
rect 298462 3176 298468 3188
rect 297416 3148 298468 3176
rect 297416 3136 297422 3148
rect 298462 3136 298468 3148
rect 298520 3136 298526 3188
rect 511350 3136 511356 3188
rect 511408 3176 511414 3188
rect 514754 3176 514760 3188
rect 511408 3148 514760 3176
rect 511408 3136 511414 3148
rect 514754 3136 514760 3148
rect 514812 3136 514818 3188
rect 122282 3068 122288 3120
rect 122340 3108 122346 3120
rect 124858 3108 124864 3120
rect 122340 3080 124864 3108
rect 122340 3068 122346 3080
rect 124858 3068 124864 3080
rect 124916 3068 124922 3120
rect 134150 3068 134156 3120
rect 134208 3108 134214 3120
rect 136818 3108 136824 3120
rect 134208 3080 136824 3108
rect 134208 3068 134214 3080
rect 136818 3068 136824 3080
rect 136876 3068 136882 3120
rect 182818 3068 182824 3120
rect 182876 3108 182882 3120
rect 184934 3108 184940 3120
rect 182876 3080 184940 3108
rect 182876 3068 182882 3080
rect 184934 3068 184940 3080
rect 184992 3068 184998 3120
rect 522298 3068 522304 3120
rect 522356 3108 522362 3120
rect 524230 3108 524236 3120
rect 522356 3080 524236 3108
rect 522356 3068 522362 3080
rect 524230 3068 524236 3080
rect 524288 3068 524294 3120
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 22738 3040 22744 3052
rect 20680 3012 22744 3040
rect 20680 3000 20686 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 23014 3000 23020 3052
rect 23072 3040 23078 3052
rect 25498 3040 25504 3052
rect 23072 3012 25504 3040
rect 23072 3000 23078 3012
rect 25498 3000 25504 3012
rect 25556 3000 25562 3052
rect 132954 3000 132960 3052
rect 133012 3040 133018 3052
rect 141418 3040 141424 3052
rect 133012 3012 141424 3040
rect 133012 3000 133018 3012
rect 141418 3000 141424 3012
rect 141476 3000 141482 3052
rect 182910 3000 182916 3052
rect 182968 3040 182974 3052
rect 189718 3040 189724 3052
rect 182968 3012 189724 3040
rect 182968 3000 182974 3012
rect 189718 3000 189724 3012
rect 189776 3000 189782 3052
rect 464338 3000 464344 3052
rect 464396 3040 464402 3052
rect 466270 3040 466276 3052
rect 464396 3012 466276 3040
rect 464396 3000 464402 3012
rect 466270 3000 466276 3012
rect 466328 3000 466334 3052
rect 514018 3000 514024 3052
rect 514076 3040 514082 3052
rect 515950 3040 515956 3052
rect 514076 3012 515956 3040
rect 514076 3000 514082 3012
rect 515950 3000 515956 3012
rect 516008 3000 516014 3052
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 14458 2972 14464 2984
rect 12400 2944 14464 2972
rect 12400 2932 12406 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 432598 2932 432604 2984
rect 432656 2972 432662 2984
rect 434438 2972 434444 2984
rect 432656 2944 434444 2972
rect 432656 2932 432662 2944
rect 434438 2932 434444 2944
rect 434496 2932 434502 2984
rect 118786 2864 118792 2916
rect 118844 2904 118850 2916
rect 122098 2904 122104 2916
rect 118844 2876 122104 2904
rect 118844 2864 118850 2876
rect 122098 2864 122104 2876
rect 122156 2864 122162 2916
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 137836 700816 137888 700868
rect 157340 700816 157392 700868
rect 155960 700748 156012 700800
rect 202788 700748 202840 700800
rect 89168 700680 89220 700732
rect 160744 700680 160796 700732
rect 154580 700612 154632 700664
rect 267648 700612 267700 700664
rect 24308 700544 24360 700596
rect 162216 700544 162268 700596
rect 8116 700476 8168 700528
rect 162124 700476 162176 700528
rect 153292 700408 153344 700460
rect 332508 700408 332560 700460
rect 152464 700340 152516 700392
rect 413652 700340 413704 700392
rect 489184 700340 489236 700392
rect 527180 700340 527232 700392
rect 527824 700340 527876 700392
rect 559656 700340 559708 700392
rect 148324 700272 148376 700324
rect 543464 700272 543516 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 396724 699660 396776 699712
rect 397460 699660 397512 699712
rect 428464 699660 428516 699712
rect 429844 699660 429896 699712
rect 146300 696940 146352 696992
rect 580172 696940 580224 696992
rect 3424 683204 3476 683256
rect 161480 683204 161532 683256
rect 146944 683136 146996 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 163504 670692 163556 670744
rect 498844 670692 498896 670744
rect 580172 670692 580224 670744
rect 3424 656888 3476 656940
rect 163596 656888 163648 656940
rect 182824 643084 182876 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 164240 632068 164292 632120
rect 188344 630640 188396 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 164884 618264 164936 618316
rect 143632 616836 143684 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 164976 605820 165028 605872
rect 142436 590656 142488 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 165620 579640 165672 579692
rect 144184 576852 144236 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 167644 565836 167696 565888
rect 142804 563048 142856 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 166264 553392 166316 553444
rect 181444 536800 181496 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 167000 527144 167052 527196
rect 142896 524424 142948 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 7564 514768 7616 514820
rect 180064 510620 180116 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 167736 500964 167788 501016
rect 139584 484372 139636 484424
rect 580172 484372 580224 484424
rect 140044 470568 140096 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 170404 462340 170456 462392
rect 178684 456764 178736 456816
rect 580172 456764 580224 456816
rect 157432 450508 157484 450560
rect 169760 450508 169812 450560
rect 3148 448536 3200 448588
rect 170496 448536 170548 448588
rect 138664 430584 138716 430636
rect 580172 430584 580224 430636
rect 3516 422288 3568 422340
rect 169760 422288 169812 422340
rect 138756 418140 138808 418192
rect 580172 418140 580224 418192
rect 2872 409844 2924 409896
rect 171784 409844 171836 409896
rect 185584 404336 185636 404388
rect 580172 404336 580224 404388
rect 3516 397468 3568 397520
rect 171876 397468 171928 397520
rect 196624 378156 196676 378208
rect 580172 378156 580224 378208
rect 2780 371288 2832 371340
rect 4804 371288 4856 371340
rect 3516 358368 3568 358420
rect 8944 358368 8996 358420
rect 135260 351908 135312 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 149704 345040 149756 345092
rect 134524 324300 134576 324352
rect 580172 324300 580224 324352
rect 3332 318792 3384 318844
rect 173900 318792 173952 318844
rect 135904 311856 135956 311908
rect 579988 311856 580040 311908
rect 3516 304988 3568 305040
rect 175924 304988 175976 305040
rect 134616 298120 134668 298172
rect 580172 298120 580224 298172
rect 3516 292544 3568 292596
rect 174544 292544 174596 292596
rect 145564 289076 145616 289128
rect 188344 289076 188396 289128
rect 149060 287648 149112 287700
rect 462320 287648 462372 287700
rect 137284 286288 137336 286340
rect 196624 286288 196676 286340
rect 150440 284928 150492 284980
rect 396724 284928 396776 284980
rect 189448 283568 189500 283620
rect 489184 283568 489236 283620
rect 147680 282888 147732 282940
rect 189080 282888 189132 282940
rect 189448 282888 189500 282940
rect 144920 282140 144972 282192
rect 182824 282140 182876 282192
rect 140780 280780 140832 280832
rect 181444 280780 181496 280832
rect 40040 279420 40092 279472
rect 160100 279420 160152 279472
rect 151084 275272 151136 275324
rect 428464 275272 428516 275324
rect 8944 273912 8996 273964
rect 173164 273912 173216 273964
rect 187700 273912 187752 273964
rect 364340 273912 364392 273964
rect 151820 273232 151872 273284
rect 187700 273232 187752 273284
rect 133144 271872 133196 271924
rect 580172 271872 580224 271924
rect 7564 271192 7616 271244
rect 169024 271192 169076 271244
rect 149152 271124 149204 271176
rect 494060 271124 494112 271176
rect 71780 269832 71832 269884
rect 158812 269832 158864 269884
rect 147772 269764 147824 269816
rect 527824 269764 527876 269816
rect 4804 268404 4856 268456
rect 172520 268404 172572 268456
rect 146208 268336 146260 268388
rect 498844 268336 498896 268388
rect 137836 266976 137888 267028
rect 185584 266976 185636 267028
rect 3056 266364 3108 266416
rect 175924 266364 175976 266416
rect 141424 265684 141476 265736
rect 180064 265684 180116 265736
rect 3424 265616 3476 265668
rect 169208 265616 169260 265668
rect 172520 265548 172572 265600
rect 190460 265548 190512 265600
rect 171876 265480 171928 265532
rect 190828 265480 190880 265532
rect 174544 265412 174596 265464
rect 194876 265412 194928 265464
rect 175832 265344 175884 265396
rect 196440 265344 196492 265396
rect 170220 265276 170272 265328
rect 170496 265276 170548 265328
rect 192024 265276 192076 265328
rect 171692 265208 171744 265260
rect 171876 265208 171928 265260
rect 173348 265208 173400 265260
rect 197636 265208 197688 265260
rect 171784 265140 171836 265192
rect 196532 265140 196584 265192
rect 169116 265072 169168 265124
rect 196256 265072 196308 265124
rect 170404 265004 170456 265056
rect 170680 265004 170732 265056
rect 197912 265004 197964 265056
rect 119712 264936 119764 264988
rect 152188 264936 152240 264988
rect 152464 264936 152516 264988
rect 160836 264936 160888 264988
rect 193404 264936 193456 264988
rect 149704 264324 149756 264376
rect 173440 264324 173492 264376
rect 139400 264256 139452 264308
rect 178684 264256 178736 264308
rect 106924 264188 106976 264240
rect 158720 264188 158772 264240
rect 119896 264052 119948 264104
rect 137836 264052 137888 264104
rect 116768 263984 116820 264036
rect 134432 263984 134484 264036
rect 134616 263984 134668 264036
rect 119528 263916 119580 263968
rect 139400 263916 139452 263968
rect 112720 263848 112772 263900
rect 133144 263848 133196 263900
rect 120908 263780 120960 263832
rect 141424 263780 141476 263832
rect 119620 263712 119672 263764
rect 142620 263712 142672 263764
rect 114008 263644 114060 263696
rect 137192 263644 137244 263696
rect 173164 263644 173216 263696
rect 173440 263644 173492 263696
rect 194968 263644 195020 263696
rect 121000 263576 121052 263628
rect 151084 263576 151136 263628
rect 158720 263576 158772 263628
rect 159364 263576 159416 263628
rect 190920 263576 190972 263628
rect 137468 263508 137520 263560
rect 580264 263508 580316 263560
rect 147680 263440 147732 263492
rect 148048 263440 148100 263492
rect 191012 263440 191064 263492
rect 282920 263440 282972 263492
rect 191840 263372 191892 263424
rect 218060 263372 218112 263424
rect 3516 263100 3568 263152
rect 176752 263100 176804 263152
rect 179236 263100 179288 263152
rect 192484 263100 192536 263152
rect 132040 263032 132092 263084
rect 580356 263032 580408 263084
rect 167828 262964 167880 263016
rect 192300 262964 192352 263016
rect 116676 262896 116728 262948
rect 127624 262896 127676 262948
rect 131120 262896 131172 262948
rect 131764 262896 131816 262948
rect 580448 262896 580500 262948
rect 3424 262828 3476 262880
rect 178408 262828 178460 262880
rect 112536 262760 112588 262812
rect 131120 262760 131172 262812
rect 166264 262760 166316 262812
rect 192208 262760 192260 262812
rect 113732 262692 113784 262744
rect 134524 262692 134576 262744
rect 134800 262692 134852 262744
rect 153200 262692 153252 262744
rect 158720 262692 158772 262744
rect 164976 262692 165028 262744
rect 193588 262692 193640 262744
rect 116584 262624 116636 262676
rect 131120 262624 131172 262676
rect 153844 262624 153896 262676
rect 188252 262624 188304 262676
rect 347780 262828 347832 262880
rect 116492 262556 116544 262608
rect 144184 262556 144236 262608
rect 155868 262556 155920 262608
rect 191012 262556 191064 262608
rect 113916 262488 113968 262540
rect 142252 262488 142304 262540
rect 142896 262488 142948 262540
rect 157156 262488 157208 262540
rect 191840 262488 191892 262540
rect 118424 262420 118476 262472
rect 125968 262420 126020 262472
rect 181812 262420 181864 262472
rect 196348 262420 196400 262472
rect 118240 262352 118292 262404
rect 129280 262352 129332 262404
rect 182916 262352 182968 262404
rect 190552 262352 190604 262404
rect 181260 262284 181312 262336
rect 190644 262284 190696 262336
rect 116860 262216 116912 262268
rect 122748 262216 122800 262268
rect 184572 262216 184624 262268
rect 189172 262216 189224 262268
rect 129832 261536 129884 261588
rect 189724 261536 189776 261588
rect 178408 261468 178460 261520
rect 200580 261468 200632 261520
rect 131120 261400 131172 261452
rect 471244 261400 471296 261452
rect 118332 261332 118384 261384
rect 127348 261332 127400 261384
rect 183468 261332 183520 261384
rect 197820 261332 197872 261384
rect 14464 261264 14516 261316
rect 176200 261264 176252 261316
rect 177304 261264 177356 261316
rect 193772 261264 193824 261316
rect 111248 261196 111300 261248
rect 134340 261196 134392 261248
rect 180524 261196 180576 261248
rect 199292 261196 199344 261248
rect 117964 261128 118016 261180
rect 127072 261128 127124 261180
rect 127348 261128 127400 261180
rect 132868 261128 132920 261180
rect 176752 261128 176804 261180
rect 196716 261128 196768 261180
rect 110880 261060 110932 261112
rect 128728 261060 128780 261112
rect 158720 261060 158772 261112
rect 193680 261060 193732 261112
rect 111064 260992 111116 261044
rect 130384 260992 130436 261044
rect 181996 260992 182048 261044
rect 200488 260992 200540 261044
rect 176200 260924 176252 260976
rect 195060 260924 195112 260976
rect 114100 260856 114152 260908
rect 125600 260856 125652 260908
rect 184020 260856 184072 260908
rect 199200 260856 199252 260908
rect 120816 260788 120868 260840
rect 123208 260788 123260 260840
rect 119804 260720 119856 260772
rect 122840 260720 122892 260772
rect 122748 260652 122800 260704
rect 124312 260652 124364 260704
rect 173900 260448 173952 260500
rect 193496 260448 193548 260500
rect 134340 260380 134392 260432
rect 188988 260380 189040 260432
rect 4804 260312 4856 260364
rect 177304 260312 177356 260364
rect 175924 260244 175976 260296
rect 192392 260244 192444 260296
rect 135260 260176 135312 260228
rect 136226 260176 136278 260228
rect 155960 260176 156012 260228
rect 156650 260176 156702 260228
rect 167000 260176 167052 260228
rect 167690 260176 167742 260228
rect 169760 260176 169812 260228
rect 171002 260176 171054 260228
rect 169208 260108 169260 260160
rect 191196 260176 191248 260228
rect 167690 260040 167742 260092
rect 189632 260040 189684 260092
rect 112628 259972 112680 260024
rect 123760 259972 123812 260024
rect 164700 259972 164752 260024
rect 189540 259972 189592 260024
rect 118148 259904 118200 259956
rect 135260 259904 135312 259956
rect 166172 259904 166224 259956
rect 191012 259904 191064 259956
rect 119344 259836 119396 259888
rect 149152 259836 149204 259888
rect 156972 259836 157024 259888
rect 189356 259836 189408 259888
rect 118056 259768 118108 259820
rect 150440 259768 150492 259820
rect 151360 259768 151412 259820
rect 171140 259768 171192 259820
rect 203248 259768 203300 259820
rect 119436 259700 119488 259752
rect 153200 259700 153252 259752
rect 158076 259700 158128 259752
rect 191104 259700 191156 259752
rect 115296 259632 115348 259684
rect 128360 259632 128412 259684
rect 184940 259632 184992 259684
rect 196624 259632 196676 259684
rect 117872 259564 117924 259616
rect 178040 259564 178092 259616
rect 195244 259564 195296 259616
rect 115480 259496 115532 259548
rect 126520 259496 126572 259548
rect 180156 259496 180208 259548
rect 197728 259496 197780 259548
rect 120724 259428 120776 259480
rect 124864 259428 124916 259480
rect 133236 259428 133288 259480
rect 472624 259428 472676 259480
rect 188988 259360 189040 259412
rect 580172 259360 580224 259412
rect 472624 245556 472676 245608
rect 580172 245556 580224 245608
rect 3516 241408 3568 241460
rect 14464 241408 14516 241460
rect 2780 215228 2832 215280
rect 4804 215228 4856 215280
rect 471244 206932 471296 206984
rect 579804 206932 579856 206984
rect 190460 200744 190512 200796
rect 128912 200676 128964 200728
rect 129280 200676 129332 200728
rect 131580 200676 131632 200728
rect 131672 200676 131724 200728
rect 178776 200676 178828 200728
rect 111616 200540 111668 200592
rect 132224 200608 132276 200660
rect 128084 200540 128136 200592
rect 131948 200540 132000 200592
rect 132040 200540 132092 200592
rect 108948 200472 109000 200524
rect 131764 200472 131816 200524
rect 130476 200404 130528 200456
rect 131856 200404 131908 200456
rect 123944 200336 123996 200388
rect 121092 200268 121144 200320
rect 131488 200200 131540 200252
rect 131764 200132 131816 200184
rect 131856 200064 131908 200116
rect 129096 199928 129148 199980
rect 132224 199928 132276 199980
rect 128360 199860 128412 199912
rect 128544 199792 128596 199844
rect 132132 199792 132184 199844
rect 131764 199724 131816 199776
rect 132546 199860 132598 199912
rect 132638 199860 132690 199912
rect 126152 199656 126204 199708
rect 133006 199860 133058 199912
rect 133190 199860 133242 199912
rect 133742 199860 133794 199912
rect 134018 199860 134070 199912
rect 134386 199860 134438 199912
rect 118516 199588 118568 199640
rect 131856 199588 131908 199640
rect 131948 199588 132000 199640
rect 133696 199724 133748 199776
rect 133972 199724 134024 199776
rect 134570 199860 134622 199912
rect 135030 199860 135082 199912
rect 135398 199860 135450 199912
rect 135582 199860 135634 199912
rect 135674 199860 135726 199912
rect 135766 199860 135818 199912
rect 134846 199792 134898 199844
rect 133144 199588 133196 199640
rect 134432 199588 134484 199640
rect 117044 199520 117096 199572
rect 131488 199520 131540 199572
rect 115664 199452 115716 199504
rect 132960 199452 133012 199504
rect 133880 199452 133932 199504
rect 134340 199452 134392 199504
rect 115756 199384 115808 199436
rect 132500 199384 132552 199436
rect 135306 199792 135358 199844
rect 134984 199588 135036 199640
rect 134800 199452 134852 199504
rect 135720 199724 135772 199776
rect 135628 199656 135680 199708
rect 136042 199860 136094 199912
rect 136226 199860 136278 199912
rect 136318 199860 136370 199912
rect 135904 199588 135956 199640
rect 136870 199860 136922 199912
rect 136962 199860 137014 199912
rect 136272 199724 136324 199776
rect 136640 199588 136692 199640
rect 135536 199520 135588 199572
rect 136548 199520 136600 199572
rect 136916 199724 136968 199776
rect 137146 199860 137198 199912
rect 137422 199860 137474 199912
rect 137514 199860 137566 199912
rect 137606 199860 137658 199912
rect 138342 199860 138394 199912
rect 138618 199860 138670 199912
rect 138710 199860 138762 199912
rect 138802 199860 138854 199912
rect 138894 199860 138946 199912
rect 137238 199792 137290 199844
rect 137100 199656 137152 199708
rect 137192 199656 137244 199708
rect 137284 199520 137336 199572
rect 137468 199724 137520 199776
rect 138848 199724 138900 199776
rect 138664 199656 138716 199708
rect 138756 199656 138808 199708
rect 139078 199792 139130 199844
rect 137652 199588 137704 199640
rect 138388 199588 138440 199640
rect 137928 199520 137980 199572
rect 139032 199520 139084 199572
rect 139216 199520 139268 199572
rect 137560 199452 137612 199504
rect 139722 199860 139774 199912
rect 139814 199860 139866 199912
rect 139906 199860 139958 199912
rect 139998 199860 140050 199912
rect 140274 199860 140326 199912
rect 140458 199860 140510 199912
rect 140734 199860 140786 199912
rect 141194 199860 141246 199912
rect 141470 199860 141522 199912
rect 139768 199656 139820 199708
rect 140044 199724 140096 199776
rect 140274 199656 140326 199708
rect 139952 199588 140004 199640
rect 140596 199588 140648 199640
rect 140780 199588 140832 199640
rect 141654 199792 141706 199844
rect 141608 199656 141660 199708
rect 141424 199588 141476 199640
rect 141838 199860 141890 199912
rect 141930 199860 141982 199912
rect 142206 199860 142258 199912
rect 141884 199724 141936 199776
rect 142160 199724 142212 199776
rect 142390 199860 142442 199912
rect 142068 199588 142120 199640
rect 142436 199588 142488 199640
rect 140780 199452 140832 199504
rect 141148 199452 141200 199504
rect 142758 199860 142810 199912
rect 143034 199860 143086 199912
rect 143126 199860 143178 199912
rect 143310 199860 143362 199912
rect 143678 199860 143730 199912
rect 143862 199860 143914 199912
rect 143954 199860 144006 199912
rect 144138 199860 144190 199912
rect 144230 199860 144282 199912
rect 142666 199792 142718 199844
rect 143218 199792 143270 199844
rect 142712 199656 142764 199708
rect 143080 199656 143132 199708
rect 143908 199724 143960 199776
rect 143264 199588 143316 199640
rect 143632 199588 143684 199640
rect 143816 199588 143868 199640
rect 144092 199588 144144 199640
rect 144184 199588 144236 199640
rect 144690 199860 144742 199912
rect 144966 199860 145018 199912
rect 145242 199860 145294 199912
rect 145702 199860 145754 199912
rect 145794 199860 145846 199912
rect 145886 199860 145938 199912
rect 145978 199860 146030 199912
rect 146070 199860 146122 199912
rect 144552 199588 144604 199640
rect 142988 199520 143040 199572
rect 145518 199792 145570 199844
rect 145610 199792 145662 199844
rect 145472 199656 145524 199708
rect 145288 199588 145340 199640
rect 145564 199588 145616 199640
rect 146116 199724 146168 199776
rect 146024 199656 146076 199708
rect 146346 199860 146398 199912
rect 146714 199860 146766 199912
rect 147174 199860 147226 199912
rect 147266 199860 147318 199912
rect 147358 199860 147410 199912
rect 147726 199860 147778 199912
rect 148094 199860 148146 199912
rect 148278 199860 148330 199912
rect 148370 199860 148422 199912
rect 145840 199588 145892 199640
rect 145932 199588 145984 199640
rect 145656 199520 145708 199572
rect 146392 199520 146444 199572
rect 146484 199520 146536 199572
rect 147220 199724 147272 199776
rect 147910 199792 147962 199844
rect 147312 199656 147364 199708
rect 147772 199656 147824 199708
rect 148048 199656 148100 199708
rect 148232 199656 148284 199708
rect 148324 199656 148376 199708
rect 148554 199860 148606 199912
rect 148554 199724 148606 199776
rect 148922 199860 148974 199912
rect 149290 199860 149342 199912
rect 149474 199860 149526 199912
rect 149566 199860 149618 199912
rect 149842 199860 149894 199912
rect 150026 199860 150078 199912
rect 150486 199860 150538 199912
rect 150578 199860 150630 199912
rect 150670 199860 150722 199912
rect 150854 199860 150906 199912
rect 150946 199860 150998 199912
rect 151038 199860 151090 199912
rect 148784 199588 148836 199640
rect 148968 199588 149020 199640
rect 149888 199724 149940 199776
rect 149520 199656 149572 199708
rect 149244 199588 149296 199640
rect 142712 199452 142764 199504
rect 144920 199452 144972 199504
rect 136456 199384 136508 199436
rect 148140 199384 148192 199436
rect 122748 199316 122800 199368
rect 130016 199316 130068 199368
rect 133144 199316 133196 199368
rect 133328 199316 133380 199368
rect 134616 199316 134668 199368
rect 139400 199316 139452 199368
rect 139768 199316 139820 199368
rect 145104 199316 145156 199368
rect 149060 199520 149112 199572
rect 149152 199520 149204 199572
rect 150302 199656 150354 199708
rect 149796 199588 149848 199640
rect 150072 199520 150124 199572
rect 150348 199520 150400 199572
rect 148968 199452 149020 199504
rect 150532 199452 150584 199504
rect 122564 199248 122616 199300
rect 145196 199248 145248 199300
rect 122472 199180 122524 199232
rect 143448 199180 143500 199232
rect 150900 199724 150952 199776
rect 151682 199860 151734 199912
rect 150808 199588 150860 199640
rect 151084 199588 151136 199640
rect 151544 199588 151596 199640
rect 150716 199384 150768 199436
rect 150900 199316 150952 199368
rect 151176 199316 151228 199368
rect 151866 199860 151918 199912
rect 151958 199860 152010 199912
rect 152326 199860 152378 199912
rect 152418 199860 152470 199912
rect 152694 199860 152746 199912
rect 152878 199860 152930 199912
rect 153154 199860 153206 199912
rect 153246 199860 153298 199912
rect 153430 199860 153482 199912
rect 153706 199860 153758 199912
rect 153890 199860 153942 199912
rect 154258 199860 154310 199912
rect 154350 199860 154402 199912
rect 155086 199860 155138 199912
rect 151912 199724 151964 199776
rect 152004 199656 152056 199708
rect 151544 199248 151596 199300
rect 152464 199656 152516 199708
rect 152970 199792 153022 199844
rect 152924 199656 152976 199708
rect 153016 199656 153068 199708
rect 152832 199520 152884 199572
rect 153660 199724 153712 199776
rect 154074 199792 154126 199844
rect 154212 199724 154264 199776
rect 153844 199588 153896 199640
rect 154028 199588 154080 199640
rect 154304 199588 154356 199640
rect 154856 199588 154908 199640
rect 155362 199860 155414 199912
rect 155316 199724 155368 199776
rect 155546 199860 155598 199912
rect 155638 199860 155690 199912
rect 156006 199860 156058 199912
rect 156098 199860 156150 199912
rect 156190 199860 156242 199912
rect 156374 199860 156426 199912
rect 156650 199860 156702 199912
rect 157386 199860 157438 199912
rect 155592 199724 155644 199776
rect 156282 199792 156334 199844
rect 156144 199724 156196 199776
rect 155868 199588 155920 199640
rect 153384 199520 153436 199572
rect 154672 199520 154724 199572
rect 155408 199520 155460 199572
rect 156052 199656 156104 199708
rect 156236 199656 156288 199708
rect 156328 199656 156380 199708
rect 157386 199724 157438 199776
rect 154856 199452 154908 199504
rect 154488 199384 154540 199436
rect 154856 199316 154908 199368
rect 156880 199384 156932 199436
rect 157156 199384 157208 199436
rect 157248 199316 157300 199368
rect 154396 199248 154448 199300
rect 154764 199248 154816 199300
rect 156972 199248 157024 199300
rect 157570 199860 157622 199912
rect 157754 199860 157806 199912
rect 157846 199860 157898 199912
rect 157938 199860 157990 199912
rect 158030 199860 158082 199912
rect 158214 199860 158266 199912
rect 158306 199860 158358 199912
rect 158490 199860 158542 199912
rect 158674 199860 158726 199912
rect 158766 199860 158818 199912
rect 158858 199860 158910 199912
rect 157800 199656 157852 199708
rect 157708 199588 157760 199640
rect 157892 199520 157944 199572
rect 158168 199588 158220 199640
rect 158444 199588 158496 199640
rect 158352 199520 158404 199572
rect 158720 199724 158772 199776
rect 158812 199724 158864 199776
rect 159134 199860 159186 199912
rect 159318 199860 159370 199912
rect 158904 199520 158956 199572
rect 178960 200404 179012 200456
rect 180248 200404 180300 200456
rect 159502 199860 159554 199912
rect 159962 199860 160014 199912
rect 160054 199860 160106 199912
rect 160146 199860 160198 199912
rect 160514 199860 160566 199912
rect 160790 199860 160842 199912
rect 160882 199860 160934 199912
rect 160974 199860 161026 199912
rect 161066 199860 161118 199912
rect 161342 199860 161394 199912
rect 161434 199860 161486 199912
rect 161710 199860 161762 199912
rect 161986 199860 162038 199912
rect 159686 199792 159738 199844
rect 159778 199792 159830 199844
rect 159870 199792 159922 199844
rect 159594 199724 159646 199776
rect 159962 199724 160014 199776
rect 159732 199656 159784 199708
rect 159824 199656 159876 199708
rect 160192 199724 160244 199776
rect 159364 199588 159416 199640
rect 159548 199588 159600 199640
rect 159180 199520 159232 199572
rect 160008 199520 160060 199572
rect 160100 199520 160152 199572
rect 160606 199792 160658 199844
rect 160836 199724 160888 199776
rect 160928 199724 160980 199776
rect 161020 199656 161072 199708
rect 161526 199792 161578 199844
rect 161388 199656 161440 199708
rect 161480 199588 161532 199640
rect 161296 199520 161348 199572
rect 161940 199656 161992 199708
rect 161848 199520 161900 199572
rect 187884 200336 187936 200388
rect 162354 199860 162406 199912
rect 162446 199860 162498 199912
rect 162538 199860 162590 199912
rect 162722 199860 162774 199912
rect 162814 199860 162866 199912
rect 162906 199860 162958 199912
rect 162676 199724 162728 199776
rect 162768 199724 162820 199776
rect 162860 199724 162912 199776
rect 162584 199588 162636 199640
rect 162400 199520 162452 199572
rect 163182 199860 163234 199912
rect 163274 199860 163326 199912
rect 163228 199656 163280 199708
rect 163320 199588 163372 199640
rect 163550 199860 163602 199912
rect 163642 199860 163694 199912
rect 163734 199860 163786 199912
rect 164010 199860 164062 199912
rect 163596 199656 163648 199708
rect 163688 199588 163740 199640
rect 163872 199588 163924 199640
rect 157984 199452 158036 199504
rect 158628 199452 158680 199504
rect 160560 199452 160612 199504
rect 160744 199452 160796 199504
rect 162308 199452 162360 199504
rect 163044 199452 163096 199504
rect 163780 199452 163832 199504
rect 159272 199384 159324 199436
rect 159640 199384 159692 199436
rect 161572 199384 161624 199436
rect 161756 199384 161808 199436
rect 162676 199384 162728 199436
rect 162860 199384 162912 199436
rect 192116 200268 192168 200320
rect 164194 199860 164246 199912
rect 164378 199792 164430 199844
rect 164516 199520 164568 199572
rect 190736 200200 190788 200252
rect 186780 200132 186832 200184
rect 164746 199860 164798 199912
rect 164930 199860 164982 199912
rect 165758 199860 165810 199912
rect 165850 199860 165902 199912
rect 165942 199860 165994 199912
rect 166126 199860 166178 199912
rect 165482 199792 165534 199844
rect 164884 199656 164936 199708
rect 165068 199588 165120 199640
rect 165804 199724 165856 199776
rect 165896 199724 165948 199776
rect 165436 199520 165488 199572
rect 164792 199452 164844 199504
rect 166494 199860 166546 199912
rect 166448 199588 166500 199640
rect 166632 199588 166684 199640
rect 166724 199588 166776 199640
rect 167046 199860 167098 199912
rect 167230 199860 167282 199912
rect 167322 199860 167374 199912
rect 167598 199860 167650 199912
rect 167966 199860 168018 199912
rect 167184 199724 167236 199776
rect 167368 199724 167420 199776
rect 167000 199588 167052 199640
rect 166356 199520 166408 199572
rect 166908 199520 166960 199572
rect 168012 199588 168064 199640
rect 166080 199452 166132 199504
rect 165620 199384 165672 199436
rect 168426 199860 168478 199912
rect 168518 199860 168570 199912
rect 168610 199860 168662 199912
rect 168794 199860 168846 199912
rect 168886 199860 168938 199912
rect 168978 199860 169030 199912
rect 169162 199860 169214 199912
rect 169254 199860 169306 199912
rect 169346 199860 169398 199912
rect 170174 199860 170226 199912
rect 170542 199860 170594 199912
rect 170634 199860 170686 199912
rect 170726 199860 170778 199912
rect 171278 199860 171330 199912
rect 171646 199860 171698 199912
rect 171738 199860 171790 199912
rect 172014 199860 172066 199912
rect 172198 199860 172250 199912
rect 168196 199520 168248 199572
rect 168564 199656 168616 199708
rect 168472 199452 168524 199504
rect 168840 199656 168892 199708
rect 168932 199656 168984 199708
rect 169208 199656 169260 199708
rect 169300 199656 169352 199708
rect 169116 199588 169168 199640
rect 170358 199792 170410 199844
rect 170588 199656 170640 199708
rect 170680 199656 170732 199708
rect 170404 199588 170456 199640
rect 170496 199588 170548 199640
rect 170864 199520 170916 199572
rect 171692 199724 171744 199776
rect 171968 199520 172020 199572
rect 172750 199860 172802 199912
rect 172842 199860 172894 199912
rect 169576 199452 169628 199504
rect 171324 199452 171376 199504
rect 172060 199452 172112 199504
rect 170036 199384 170088 199436
rect 171876 199384 171928 199436
rect 173026 199860 173078 199912
rect 178500 200064 178552 200116
rect 173302 199860 173354 199912
rect 173578 199860 173630 199912
rect 173854 199860 173906 199912
rect 173946 199860 173998 199912
rect 174590 199860 174642 199912
rect 174682 199860 174734 199912
rect 172980 199520 173032 199572
rect 172428 199452 172480 199504
rect 172796 199452 172848 199504
rect 172888 199384 172940 199436
rect 174130 199792 174182 199844
rect 173992 199588 174044 199640
rect 174176 199588 174228 199640
rect 173808 199520 173860 199572
rect 173900 199520 173952 199572
rect 173440 199452 173492 199504
rect 173716 199452 173768 199504
rect 174636 199656 174688 199708
rect 178132 199996 178184 200048
rect 174958 199860 175010 199912
rect 175142 199860 175194 199912
rect 175326 199860 175378 199912
rect 174820 199588 174872 199640
rect 175280 199588 175332 199640
rect 177948 199928 178000 199980
rect 175510 199860 175562 199912
rect 176062 199860 176114 199912
rect 176246 199860 176298 199912
rect 176430 199860 176482 199912
rect 176706 199860 176758 199912
rect 176890 199860 176942 199912
rect 176982 199860 177034 199912
rect 177074 199860 177126 199912
rect 175096 199520 175148 199572
rect 175004 199452 175056 199504
rect 176200 199588 176252 199640
rect 176660 199656 176712 199708
rect 176476 199588 176528 199640
rect 177028 199724 177080 199776
rect 176936 199656 176988 199708
rect 176844 199520 176896 199572
rect 177304 199520 177356 199572
rect 188160 199520 188212 199572
rect 177672 199452 177724 199504
rect 182916 199452 182968 199504
rect 190552 199452 190604 199504
rect 179328 199384 179380 199436
rect 180892 199384 180944 199436
rect 190644 199384 190696 199436
rect 167644 199316 167696 199368
rect 170312 199316 170364 199368
rect 200396 199316 200448 199368
rect 164792 199248 164844 199300
rect 167368 199248 167420 199300
rect 201684 199248 201736 199300
rect 155316 199180 155368 199232
rect 160008 199180 160060 199232
rect 170404 199180 170456 199232
rect 172152 199180 172204 199232
rect 180156 199180 180208 199232
rect 180800 199180 180852 199232
rect 189816 199180 189868 199232
rect 122380 199112 122432 199164
rect 145656 199112 145708 199164
rect 155868 199112 155920 199164
rect 189080 199112 189132 199164
rect 121184 199044 121236 199096
rect 132776 199044 132828 199096
rect 132960 199044 133012 199096
rect 147588 199044 147640 199096
rect 150992 199044 151044 199096
rect 158536 199044 158588 199096
rect 121276 198976 121328 199028
rect 146576 198976 146628 199028
rect 153660 198976 153712 199028
rect 162308 199044 162360 199096
rect 163136 199044 163188 199096
rect 197544 199044 197596 199096
rect 158996 198976 159048 199028
rect 193220 198976 193272 199028
rect 129556 198908 129608 198960
rect 139032 198908 139084 198960
rect 139952 198908 140004 198960
rect 144184 198908 144236 198960
rect 153936 198908 153988 198960
rect 187792 198908 187844 198960
rect 129188 198840 129240 198892
rect 147956 198840 148008 198892
rect 165988 198840 166040 198892
rect 166724 198840 166776 198892
rect 126336 198772 126388 198824
rect 144552 198772 144604 198824
rect 157248 198772 157300 198824
rect 166080 198772 166132 198824
rect 170312 198840 170364 198892
rect 170404 198840 170456 198892
rect 172152 198840 172204 198892
rect 169760 198772 169812 198824
rect 174452 198840 174504 198892
rect 172428 198772 172480 198824
rect 172980 198772 173032 198824
rect 173256 198772 173308 198824
rect 174820 198840 174872 198892
rect 175464 198840 175516 198892
rect 180800 198840 180852 198892
rect 174636 198772 174688 198824
rect 175648 198772 175700 198824
rect 175740 198772 175792 198824
rect 176752 198772 176804 198824
rect 177948 198772 178000 198824
rect 187516 198840 187568 198892
rect 183836 198772 183888 198824
rect 189172 198772 189224 198824
rect 122656 198704 122708 198756
rect 135076 198636 135128 198688
rect 135260 198636 135312 198688
rect 143724 198704 143776 198756
rect 144092 198704 144144 198756
rect 166632 198704 166684 198756
rect 171416 198704 171468 198756
rect 146208 198636 146260 198688
rect 167184 198636 167236 198688
rect 174176 198636 174228 198688
rect 175924 198704 175976 198756
rect 176476 198704 176528 198756
rect 177672 198704 177724 198756
rect 201040 198704 201092 198756
rect 188344 198636 188396 198688
rect 123116 198568 123168 198620
rect 143632 198568 143684 198620
rect 148508 198568 148560 198620
rect 149428 198568 149480 198620
rect 156788 198568 156840 198620
rect 157156 198568 157208 198620
rect 167092 198568 167144 198620
rect 170496 198568 170548 198620
rect 171876 198568 171928 198620
rect 187056 198568 187108 198620
rect 108580 198500 108632 198552
rect 129004 198500 129056 198552
rect 131764 198500 131816 198552
rect 137560 198500 137612 198552
rect 137744 198500 137796 198552
rect 138020 198500 138072 198552
rect 145656 198500 145708 198552
rect 156696 198500 156748 198552
rect 171140 198500 171192 198552
rect 186872 198500 186924 198552
rect 131856 198432 131908 198484
rect 107108 198364 107160 198416
rect 128544 198364 128596 198416
rect 130384 198364 130436 198416
rect 138940 198364 138992 198416
rect 141516 198432 141568 198484
rect 142068 198432 142120 198484
rect 157800 198432 157852 198484
rect 172428 198432 172480 198484
rect 174176 198432 174228 198484
rect 178316 198432 178368 198484
rect 147680 198364 147732 198416
rect 157064 198364 157116 198416
rect 157432 198364 157484 198416
rect 158076 198364 158128 198416
rect 173440 198364 173492 198416
rect 108672 198296 108724 198348
rect 136456 198296 136508 198348
rect 136548 198296 136600 198348
rect 145840 198296 145892 198348
rect 156420 198296 156472 198348
rect 122104 198228 122156 198280
rect 148508 198228 148560 198280
rect 151728 198228 151780 198280
rect 158720 198228 158772 198280
rect 170220 198296 170272 198348
rect 187976 198364 188028 198416
rect 174452 198296 174504 198348
rect 186964 198296 187016 198348
rect 104440 198160 104492 198212
rect 133236 198160 133288 198212
rect 138020 198160 138072 198212
rect 139860 198160 139912 198212
rect 103060 198092 103112 198144
rect 133972 198092 134024 198144
rect 103152 198024 103204 198076
rect 128912 198024 128964 198076
rect 132776 198024 132828 198076
rect 146024 198092 146076 198144
rect 170772 198228 170824 198280
rect 188068 198228 188120 198280
rect 170404 198160 170456 198212
rect 188436 198160 188488 198212
rect 140780 198024 140832 198076
rect 141148 198024 141200 198076
rect 155960 198024 156012 198076
rect 171048 198092 171100 198144
rect 172520 198092 172572 198144
rect 172704 198092 172756 198144
rect 173900 198092 173952 198144
rect 195336 198092 195388 198144
rect 171140 198024 171192 198076
rect 171324 198024 171376 198076
rect 173256 198024 173308 198076
rect 102784 197956 102836 198008
rect 126152 197956 126204 198008
rect 139492 197956 139544 198008
rect 140504 197956 140556 198008
rect 165344 197956 165396 198008
rect 174176 197956 174228 198008
rect 175648 197956 175700 198008
rect 198096 198024 198148 198076
rect 178500 197956 178552 198008
rect 199108 197956 199160 198008
rect 128268 197888 128320 197940
rect 148048 197888 148100 197940
rect 155408 197888 155460 197940
rect 171600 197888 171652 197940
rect 179328 197888 179380 197940
rect 186688 197888 186740 197940
rect 132224 197820 132276 197872
rect 151452 197820 151504 197872
rect 173808 197820 173860 197872
rect 187424 197820 187476 197872
rect 126796 197752 126848 197804
rect 145288 197752 145340 197804
rect 159640 197752 159692 197804
rect 173716 197752 173768 197804
rect 126704 197684 126756 197736
rect 146668 197684 146720 197736
rect 153384 197684 153436 197736
rect 179052 197684 179104 197736
rect 123668 197616 123720 197668
rect 145104 197616 145156 197668
rect 165436 197616 165488 197668
rect 178960 197616 179012 197668
rect 132776 197548 132828 197600
rect 145932 197548 145984 197600
rect 175280 197548 175332 197600
rect 175556 197548 175608 197600
rect 134800 197480 134852 197532
rect 135352 197480 135404 197532
rect 136640 197480 136692 197532
rect 137192 197480 137244 197532
rect 161480 197480 161532 197532
rect 161756 197480 161808 197532
rect 167736 197480 167788 197532
rect 180616 197480 180668 197532
rect 162676 197412 162728 197464
rect 163044 197412 163096 197464
rect 144552 197344 144604 197396
rect 146944 197344 146996 197396
rect 147036 197344 147088 197396
rect 147312 197344 147364 197396
rect 161480 197344 161532 197396
rect 162032 197344 162084 197396
rect 162952 197344 163004 197396
rect 163320 197344 163372 197396
rect 165712 197344 165764 197396
rect 165988 197344 166040 197396
rect 171232 197344 171284 197396
rect 171416 197344 171468 197396
rect 174084 197344 174136 197396
rect 174360 197344 174412 197396
rect 175280 197344 175332 197396
rect 175832 197344 175884 197396
rect 113824 197276 113876 197328
rect 139216 197276 139268 197328
rect 160100 197276 160152 197328
rect 161204 197276 161256 197328
rect 175372 197276 175424 197328
rect 176568 197276 176620 197328
rect 176660 197276 176712 197328
rect 179144 197276 179196 197328
rect 114192 197208 114244 197260
rect 143172 197208 143224 197260
rect 163964 197208 164016 197260
rect 194692 197208 194744 197260
rect 108396 197140 108448 197192
rect 132960 197140 133012 197192
rect 114468 197072 114520 197124
rect 132776 197072 132828 197124
rect 107200 197004 107252 197056
rect 138296 197140 138348 197192
rect 162216 197140 162268 197192
rect 194784 197140 194836 197192
rect 163504 197072 163556 197124
rect 197360 197072 197412 197124
rect 133236 197004 133288 197056
rect 144000 197004 144052 197056
rect 162860 197004 162912 197056
rect 163780 197004 163832 197056
rect 168472 197004 168524 197056
rect 168840 197004 168892 197056
rect 178960 197004 179012 197056
rect 198832 197004 198884 197056
rect 111156 196936 111208 196988
rect 142252 196936 142304 196988
rect 161940 196936 161992 196988
rect 196072 196936 196124 196988
rect 117136 196868 117188 196920
rect 149980 196868 150032 196920
rect 163872 196868 163924 196920
rect 197452 196868 197504 196920
rect 110236 196800 110288 196852
rect 144276 196800 144328 196852
rect 161388 196800 161440 196852
rect 194600 196800 194652 196852
rect 106004 196732 106056 196784
rect 139676 196732 139728 196784
rect 174176 196732 174228 196784
rect 199016 196732 199068 196784
rect 110052 196664 110104 196716
rect 133144 196664 133196 196716
rect 161664 196664 161716 196716
rect 162400 196664 162452 196716
rect 164424 196664 164476 196716
rect 198924 196664 198976 196716
rect 109960 196596 110012 196648
rect 133236 196596 133288 196648
rect 161848 196596 161900 196648
rect 196164 196596 196216 196648
rect 124864 196528 124916 196580
rect 151084 196528 151136 196580
rect 123024 196460 123076 196512
rect 143356 196460 143408 196512
rect 172428 196460 172480 196512
rect 191932 196460 191984 196512
rect 129280 196392 129332 196444
rect 145472 196392 145524 196444
rect 160008 196392 160060 196444
rect 169944 196392 169996 196444
rect 173440 196392 173492 196444
rect 191840 196392 191892 196444
rect 133144 196324 133196 196376
rect 144644 196324 144696 196376
rect 164516 196324 164568 196376
rect 180524 196324 180576 196376
rect 132960 196256 133012 196308
rect 137744 196256 137796 196308
rect 160376 196256 160428 196308
rect 169760 196256 169812 196308
rect 161112 196188 161164 196240
rect 182824 196188 182876 196240
rect 160836 196120 160888 196172
rect 183192 196120 183244 196172
rect 160376 196052 160428 196104
rect 160928 196052 160980 196104
rect 171140 196052 171192 196104
rect 171876 196052 171928 196104
rect 128728 195984 128780 196036
rect 142436 195984 142488 196036
rect 146760 195984 146812 196036
rect 147404 195984 147456 196036
rect 162768 195984 162820 196036
rect 167000 195984 167052 196036
rect 112996 195916 113048 195968
rect 142896 195916 142948 195968
rect 158904 195916 158956 195968
rect 159824 195916 159876 195968
rect 171048 195916 171100 195968
rect 190644 195916 190696 195968
rect 112812 195848 112864 195900
rect 143080 195848 143132 195900
rect 156052 195848 156104 195900
rect 157156 195848 157208 195900
rect 171876 195848 171928 195900
rect 172152 195848 172204 195900
rect 172612 195848 172664 195900
rect 172888 195848 172940 195900
rect 173716 195848 173768 195900
rect 193312 195848 193364 195900
rect 108764 195780 108816 195832
rect 140688 195780 140740 195832
rect 165620 195780 165672 195832
rect 183284 195780 183336 195832
rect 108488 195712 108540 195764
rect 140504 195712 140556 195764
rect 162676 195712 162728 195764
rect 183008 195712 183060 195764
rect 100668 195644 100720 195696
rect 133328 195644 133380 195696
rect 133972 195644 134024 195696
rect 141056 195644 141108 195696
rect 159088 195644 159140 195696
rect 159548 195644 159600 195696
rect 111524 195576 111576 195628
rect 144092 195576 144144 195628
rect 154212 195576 154264 195628
rect 112904 195508 112956 195560
rect 145012 195508 145064 195560
rect 158628 195508 158680 195560
rect 180248 195644 180300 195696
rect 172060 195576 172112 195628
rect 195152 195576 195204 195628
rect 101680 195440 101732 195492
rect 134156 195440 134208 195492
rect 172152 195508 172204 195560
rect 177304 195508 177356 195560
rect 190460 195440 190512 195492
rect 105728 195372 105780 195424
rect 139308 195372 139360 195424
rect 156604 195372 156656 195424
rect 131856 195304 131908 195356
rect 133972 195304 134024 195356
rect 134064 195304 134116 195356
rect 134984 195304 135036 195356
rect 152924 195304 152976 195356
rect 121368 195236 121420 195288
rect 132040 195236 132092 195288
rect 134248 195236 134300 195288
rect 134616 195236 134668 195288
rect 158076 195236 158128 195288
rect 158444 195236 158496 195288
rect 158812 195304 158864 195356
rect 159364 195304 159416 195356
rect 162584 195372 162636 195424
rect 195980 195372 196032 195424
rect 190552 195304 190604 195356
rect 186596 195236 186648 195288
rect 122196 195168 122248 195220
rect 148324 195168 148376 195220
rect 165620 195168 165672 195220
rect 166724 195168 166776 195220
rect 169760 195168 169812 195220
rect 172060 195168 172112 195220
rect 176844 195168 176896 195220
rect 177212 195168 177264 195220
rect 177304 195168 177356 195220
rect 189264 195168 189316 195220
rect 122288 195100 122340 195152
rect 144828 195100 144880 195152
rect 164424 195100 164476 195152
rect 165160 195100 165212 195152
rect 176752 195100 176804 195152
rect 177580 195100 177632 195152
rect 126428 195032 126480 195084
rect 144092 195032 144144 195084
rect 176660 195032 176712 195084
rect 177672 195032 177724 195084
rect 121920 194964 121972 195016
rect 156788 194964 156840 195016
rect 165712 194964 165764 195016
rect 166448 194964 166500 195016
rect 171508 194964 171560 195016
rect 189172 194964 189224 195016
rect 156144 194896 156196 194948
rect 180432 194896 180484 194948
rect 106188 194488 106240 194540
rect 136732 194488 136784 194540
rect 105912 194420 105964 194472
rect 136916 194420 136968 194472
rect 103244 194352 103296 194404
rect 135168 194352 135220 194404
rect 104532 194284 104584 194336
rect 136088 194284 136140 194336
rect 104624 194216 104676 194268
rect 135444 194216 135496 194268
rect 104164 194148 104216 194200
rect 135904 194148 135956 194200
rect 102968 194080 103020 194132
rect 134892 194080 134944 194132
rect 107016 194012 107068 194064
rect 138020 194012 138072 194064
rect 103428 193944 103480 193996
rect 136364 193944 136416 193996
rect 103336 193876 103388 193928
rect 136640 193876 136692 193928
rect 168840 193876 168892 193928
rect 203156 193876 203208 193928
rect 105820 193808 105872 193860
rect 140228 193808 140280 193860
rect 168196 193808 168248 193860
rect 201868 193808 201920 193860
rect 106924 193740 106976 193792
rect 137468 193740 137520 193792
rect 104072 193672 104124 193724
rect 128360 193672 128412 193724
rect 123392 193604 123444 193656
rect 148232 193604 148284 193656
rect 145564 193196 145616 193248
rect 149612 193196 149664 193248
rect 127716 193128 127768 193180
rect 139492 193128 139544 193180
rect 163320 193128 163372 193180
rect 179236 193128 179288 193180
rect 189724 193128 189776 193180
rect 580172 193128 580224 193180
rect 114376 193060 114428 193112
rect 144000 193060 144052 193112
rect 154396 193060 154448 193112
rect 181536 193060 181588 193112
rect 115388 192992 115440 193044
rect 146116 192992 146168 193044
rect 153292 192992 153344 193044
rect 181628 192992 181680 193044
rect 101864 192924 101916 192976
rect 134708 192924 134760 192976
rect 165436 192924 165488 192976
rect 193864 192924 193916 192976
rect 116952 192856 117004 192908
rect 149612 192856 149664 192908
rect 172888 192856 172940 192908
rect 206100 192856 206152 192908
rect 111432 192788 111484 192840
rect 143908 192788 143960 192840
rect 169392 192788 169444 192840
rect 202880 192788 202932 192840
rect 109776 192720 109828 192772
rect 142620 192720 142672 192772
rect 169024 192720 169076 192772
rect 203064 192720 203116 192772
rect 117228 192652 117280 192704
rect 150532 192652 150584 192704
rect 179696 192652 179748 192704
rect 202420 192652 202472 192704
rect 108856 192584 108908 192636
rect 142068 192584 142120 192636
rect 168748 192584 168800 192636
rect 202972 192584 203024 192636
rect 109868 192516 109920 192568
rect 144184 192516 144236 192568
rect 156328 192516 156380 192568
rect 205640 192516 205692 192568
rect 112444 192448 112496 192500
rect 144552 192448 144604 192500
rect 150716 192448 150768 192500
rect 206192 192448 206244 192500
rect 114836 192380 114888 192432
rect 144644 192380 144696 192432
rect 170496 192380 170548 192432
rect 196808 192380 196860 192432
rect 127808 192312 127860 192364
rect 139860 192312 139912 192364
rect 180616 192312 180668 192364
rect 201592 192312 201644 192364
rect 130568 192244 130620 192296
rect 140044 192244 140096 192296
rect 165804 192244 165856 192296
rect 178960 192244 179012 192296
rect 149704 192176 149756 192228
rect 151820 192176 151872 192228
rect 148968 191496 149020 191548
rect 157616 191496 157668 191548
rect 115572 191428 115624 191480
rect 139124 191428 139176 191480
rect 113088 191360 113140 191412
rect 138940 191360 138992 191412
rect 111708 191292 111760 191344
rect 138112 191292 138164 191344
rect 110328 191224 110380 191276
rect 138388 191224 138440 191276
rect 150624 191224 150676 191276
rect 151544 191224 151596 191276
rect 167276 191224 167328 191276
rect 168288 191224 168340 191276
rect 104808 191156 104860 191208
rect 137652 191156 137704 191208
rect 153292 191156 153344 191208
rect 154304 191156 154356 191208
rect 169944 191156 169996 191208
rect 170864 191156 170916 191208
rect 172520 191156 172572 191208
rect 173348 191156 173400 191208
rect 174084 191156 174136 191208
rect 174728 191156 174780 191208
rect 104348 191088 104400 191140
rect 138664 191088 138716 191140
rect 169852 191088 169904 191140
rect 170588 191088 170640 191140
rect 171324 191088 171376 191140
rect 171968 191088 172020 191140
rect 172704 191088 172756 191140
rect 173624 191088 173676 191140
rect 173992 191088 174044 191140
rect 174452 191088 174504 191140
rect 175372 191088 175424 191140
rect 176108 191088 176160 191140
rect 135628 191020 135680 191072
rect 136180 191020 136232 191072
rect 142620 191020 142672 191072
rect 143264 191020 143316 191072
rect 168472 191020 168524 191072
rect 169208 191020 169260 191072
rect 170036 191020 170088 191072
rect 170220 191020 170272 191072
rect 173900 191020 173952 191072
rect 175004 191020 175056 191072
rect 110144 190136 110196 190188
rect 141700 190136 141752 190188
rect 102876 190068 102928 190120
rect 135536 190068 135588 190120
rect 101588 190000 101640 190052
rect 134064 190000 134116 190052
rect 164332 190000 164384 190052
rect 164608 190000 164660 190052
rect 108120 189932 108172 189984
rect 141240 189932 141292 189984
rect 101956 189864 102008 189916
rect 135812 189864 135864 189916
rect 171232 189864 171284 189916
rect 172244 189864 172296 189916
rect 101772 189796 101824 189848
rect 135352 189796 135404 189848
rect 106832 189728 106884 189780
rect 141884 189728 141936 189780
rect 147588 189116 147640 189168
rect 154764 189116 154816 189168
rect 3424 188980 3476 189032
rect 117872 188980 117924 189032
rect 154856 187552 154908 187604
rect 155684 187552 155736 187604
rect 160560 186872 160612 186924
rect 180064 186872 180116 186924
rect 148600 185784 148652 185836
rect 154672 185784 154724 185836
rect 152556 185648 152608 185700
rect 153016 185648 153068 185700
rect 154764 185580 154816 185632
rect 155500 185580 155552 185632
rect 153384 185444 153436 185496
rect 154120 185444 154172 185496
rect 160192 185376 160244 185428
rect 160652 185376 160704 185428
rect 148048 184900 148100 184952
rect 148876 184900 148928 184952
rect 145748 184696 145800 184748
rect 156236 184696 156288 184748
rect 126612 183472 126664 183524
rect 137928 183472 137980 183524
rect 149796 183200 149848 183252
rect 151176 183200 151228 183252
rect 163136 182384 163188 182436
rect 163688 182384 163740 182436
rect 188528 178032 188580 178084
rect 580172 178032 580224 178084
rect 189724 165588 189776 165640
rect 580172 165588 580224 165640
rect 193772 156612 193824 156664
rect 193956 156612 194008 156664
rect 168564 155388 168616 155440
rect 203340 155388 203392 155440
rect 168656 155320 168708 155372
rect 203524 155320 203576 155372
rect 168472 155252 168524 155304
rect 203432 155252 203484 155304
rect 167276 155184 167328 155236
rect 202328 155184 202380 155236
rect 161756 153144 161808 153196
rect 184664 153144 184716 153196
rect 160468 153076 160520 153128
rect 184204 153076 184256 153128
rect 161572 153008 161624 153060
rect 185584 153008 185636 153060
rect 160376 152940 160428 152992
rect 185768 152940 185820 152992
rect 163044 152872 163096 152924
rect 198188 152872 198240 152924
rect 164516 152804 164568 152856
rect 199568 152804 199620 152856
rect 165988 152736 166040 152788
rect 200672 152736 200724 152788
rect 168380 152668 168432 152720
rect 203800 152668 203852 152720
rect 167092 152600 167144 152652
rect 202052 152600 202104 152652
rect 168288 152532 168340 152584
rect 202236 152532 202288 152584
rect 162768 152464 162820 152516
rect 202144 152464 202196 152516
rect 163228 152396 163280 152448
rect 184296 152396 184348 152448
rect 160284 150356 160336 150408
rect 185768 150356 185820 150408
rect 158996 150288 159048 150340
rect 184388 150288 184440 150340
rect 158904 150220 158956 150272
rect 184572 150220 184624 150272
rect 158812 150152 158864 150204
rect 184756 150152 184808 150204
rect 176844 150084 176896 150136
rect 203708 150084 203760 150136
rect 176936 150016 176988 150068
rect 204352 150016 204404 150068
rect 175648 149948 175700 150000
rect 203616 149948 203668 150000
rect 175464 149880 175516 149932
rect 204536 149880 204588 149932
rect 171600 149812 171652 149864
rect 203248 149812 203300 149864
rect 152096 149744 152148 149796
rect 204628 149744 204680 149796
rect 149244 149676 149296 149728
rect 204444 149676 204496 149728
rect 159088 149608 159140 149660
rect 184480 149608 184532 149660
rect 3424 149064 3476 149116
rect 9588 149064 9640 149116
rect 115020 148996 115072 149048
rect 142620 148996 142672 149048
rect 165620 148996 165672 149048
rect 187148 148996 187200 149048
rect 113548 148928 113600 148980
rect 143080 148928 143132 148980
rect 161480 148928 161532 148980
rect 195428 148928 195480 148980
rect 125048 148860 125100 148912
rect 153384 148860 153436 148912
rect 165896 148860 165948 148912
rect 200948 148860 201000 148912
rect 120448 148792 120500 148844
rect 149796 148792 149848 148844
rect 166908 148792 166960 148844
rect 200856 148792 200908 148844
rect 108212 148724 108264 148776
rect 138388 148724 138440 148776
rect 164424 148724 164476 148776
rect 199660 148724 199712 148776
rect 122012 148656 122064 148708
rect 153476 148656 153528 148708
rect 167828 148656 167880 148708
rect 201960 148656 202012 148708
rect 100208 148588 100260 148640
rect 133696 148588 133748 148640
rect 162952 148588 163004 148640
rect 198464 148588 198516 148640
rect 100392 148520 100444 148572
rect 134248 148520 134300 148572
rect 165712 148520 165764 148572
rect 200764 148520 200816 148572
rect 100300 148452 100352 148504
rect 134432 148452 134484 148504
rect 164332 148452 164384 148504
rect 199476 148452 199528 148504
rect 105636 148384 105688 148436
rect 139768 148384 139820 148436
rect 164240 148384 164292 148436
rect 199384 148384 199436 148436
rect 9588 148316 9640 148368
rect 180892 148316 180944 148368
rect 199292 148316 199344 148368
rect 121736 148248 121788 148300
rect 148324 148248 148376 148300
rect 179236 148248 179288 148300
rect 194140 148248 194192 148300
rect 114928 148180 114980 148232
rect 140964 148180 141016 148232
rect 112260 148112 112312 148164
rect 135628 148112 135680 148164
rect 179144 147568 179196 147620
rect 196440 147568 196492 147620
rect 171508 147500 171560 147552
rect 179236 147500 179288 147552
rect 179328 147500 179380 147552
rect 196532 147500 196584 147552
rect 178408 147432 178460 147484
rect 197912 147432 197964 147484
rect 170128 147364 170180 147416
rect 192760 147364 192812 147416
rect 178224 147296 178276 147348
rect 200580 147296 200632 147348
rect 117964 147228 118016 147280
rect 127532 147228 127584 147280
rect 115204 147160 115256 147212
rect 131856 147160 131908 147212
rect 110880 147092 110932 147144
rect 128360 147092 128412 147144
rect 117688 147024 117740 147076
rect 142528 147024 142580 147076
rect 110880 146956 110932 147008
rect 137100 146956 137152 147008
rect 117596 146888 117648 146940
rect 146484 146888 146536 146940
rect 148600 146888 148652 146940
rect 178684 147228 178736 147280
rect 179236 147228 179288 147280
rect 194048 147228 194100 147280
rect 172980 147160 173032 147212
rect 178776 147160 178828 147212
rect 172612 147092 172664 147144
rect 196992 147160 197044 147212
rect 179236 147092 179288 147144
rect 195520 147092 195572 147144
rect 172888 147024 172940 147076
rect 197084 147024 197136 147076
rect 178868 146956 178920 147008
rect 179052 146956 179104 147008
rect 172796 146820 172848 146872
rect 198280 146956 198332 147008
rect 171416 146752 171468 146804
rect 179236 146752 179288 146804
rect 178040 146684 178092 146736
rect 196716 146888 196768 146940
rect 180524 146820 180576 146872
rect 192852 146820 192904 146872
rect 128360 146344 128412 146396
rect 580448 146344 580500 146396
rect 127532 146276 127584 146328
rect 580264 146276 580316 146328
rect 113456 146208 113508 146260
rect 127808 146208 127860 146260
rect 179512 146208 179564 146260
rect 195060 146208 195112 146260
rect 115296 146140 115348 146192
rect 128912 146140 128964 146192
rect 183836 146140 183888 146192
rect 199200 146140 199252 146192
rect 112720 146072 112772 146124
rect 129924 146072 129976 146124
rect 178316 146072 178368 146124
rect 193956 146072 194008 146124
rect 112536 146004 112588 146056
rect 131304 146004 131356 146056
rect 178592 146004 178644 146056
rect 195244 146004 195296 146056
rect 113732 145936 113784 145988
rect 131580 145936 131632 145988
rect 175280 145936 175332 145988
rect 195336 145936 195388 145988
rect 112536 145868 112588 145920
rect 131764 145868 131816 145920
rect 172520 145868 172572 145920
rect 195060 145868 195112 145920
rect 119068 145800 119120 145852
rect 151452 145800 151504 145852
rect 173992 145800 174044 145852
rect 198004 145800 198056 145852
rect 117504 145732 117556 145784
rect 149704 145732 149756 145784
rect 160192 145732 160244 145784
rect 192944 145732 192996 145784
rect 118976 145664 119028 145716
rect 153016 145664 153068 145716
rect 160652 145664 160704 145716
rect 193404 145664 193456 145716
rect 116216 145596 116268 145648
rect 147864 145596 147916 145648
rect 148968 145596 149020 145648
rect 190000 145596 190052 145648
rect 3516 145528 3568 145580
rect 183468 145528 183520 145580
rect 200488 145528 200540 145580
rect 179420 145460 179472 145512
rect 194876 145460 194928 145512
rect 179604 145392 179656 145444
rect 192484 145392 192536 145444
rect 120540 144916 120592 144968
rect 182272 144916 182324 144968
rect 183468 144916 183520 144968
rect 184664 144848 184716 144900
rect 196900 144848 196952 144900
rect 172428 144780 172480 144832
rect 190828 144780 190880 144832
rect 112720 144712 112772 144764
rect 130384 144712 130436 144764
rect 173808 144712 173860 144764
rect 194968 144712 195020 144764
rect 110788 144644 110840 144696
rect 130568 144644 130620 144696
rect 169668 144644 169720 144696
rect 196256 144644 196308 144696
rect 114008 144576 114060 144628
rect 137008 144576 137060 144628
rect 165528 144576 165580 144628
rect 193588 144576 193640 144628
rect 116492 144508 116544 144560
rect 144184 144508 144236 144560
rect 160100 144508 160152 144560
rect 194232 144508 194284 144560
rect 113916 144440 113968 144492
rect 142528 144440 142580 144492
rect 162492 144440 162544 144492
rect 193404 144440 193456 144492
rect 119712 144372 119764 144424
rect 152464 144372 152516 144424
rect 159456 144372 159508 144424
rect 193680 144372 193732 144424
rect 117872 144304 117924 144356
rect 151912 144304 151964 144356
rect 154488 144304 154540 144356
rect 188252 144304 188304 144356
rect 111064 144236 111116 144288
rect 131212 144236 131264 144288
rect 188528 144236 188580 144288
rect 118240 144168 118292 144220
rect 130200 144168 130252 144220
rect 189724 144168 189776 144220
rect 180340 144100 180392 144152
rect 191288 144100 191340 144152
rect 118332 143556 118384 143608
rect 145288 143556 145340 143608
rect 116676 143488 116728 143540
rect 128452 143488 128504 143540
rect 128912 143488 128964 143540
rect 580356 143488 580408 143540
rect 114008 143420 114060 143472
rect 127716 143420 127768 143472
rect 129740 143420 129792 143472
rect 137560 143420 137612 143472
rect 146300 143420 146352 143472
rect 149152 143420 149204 143472
rect 176292 143420 176344 143472
rect 179144 143420 179196 143472
rect 180432 143420 180484 143472
rect 191472 143420 191524 143472
rect 118424 143352 118476 143404
rect 133144 143352 133196 143404
rect 172888 143352 172940 143404
rect 179328 143352 179380 143404
rect 185676 143352 185728 143404
rect 196624 143352 196676 143404
rect 116584 143284 116636 143336
rect 131488 143284 131540 143336
rect 131580 143284 131632 143336
rect 135444 143284 135496 143336
rect 171048 143284 171100 143336
rect 178408 143284 178460 143336
rect 181536 143284 181588 143336
rect 190092 143284 190144 143336
rect 190184 143284 190236 143336
rect 198372 143284 198424 143336
rect 116768 143216 116820 143268
rect 134800 143216 134852 143268
rect 175740 143216 175792 143268
rect 179420 143216 179472 143268
rect 183744 143216 183796 143268
rect 197820 143216 197872 143268
rect 118148 143148 118200 143200
rect 136640 143148 136692 143200
rect 176568 143148 176620 143200
rect 192392 143148 192444 143200
rect 120908 143080 120960 143132
rect 141608 143080 141660 143132
rect 170220 143080 170272 143132
rect 191196 143080 191248 143132
rect 119528 143012 119580 143064
rect 139768 143012 139820 143064
rect 168288 143012 168340 143064
rect 184112 143012 184164 143064
rect 184296 143012 184348 143064
rect 190184 143012 190236 143064
rect 119620 142944 119672 142996
rect 143080 142944 143132 142996
rect 174636 142944 174688 142996
rect 197636 142944 197688 142996
rect 111248 142876 111300 142928
rect 134248 142876 134300 142928
rect 166908 142876 166960 142928
rect 191012 142876 191064 142928
rect 108120 142808 108172 142860
rect 116492 142808 116544 142860
rect 121000 142808 121052 142860
rect 151360 142808 151412 142860
rect 158628 142808 158680 142860
rect 191104 142808 191156 142860
rect 118332 142740 118384 142792
rect 112628 142672 112680 142724
rect 124312 142672 124364 142724
rect 129832 142740 129884 142792
rect 135904 142740 135956 142792
rect 178132 142740 178184 142792
rect 178592 142740 178644 142792
rect 184112 142740 184164 142792
rect 189632 142740 189684 142792
rect 130476 142672 130528 142724
rect 177396 142672 177448 142724
rect 179512 142672 179564 142724
rect 178224 142536 178276 142588
rect 187700 142536 187752 142588
rect 129924 142196 129976 142248
rect 133880 142196 133932 142248
rect 155592 142196 155644 142248
rect 157340 142196 157392 142248
rect 159180 142196 159232 142248
rect 161480 142196 161532 142248
rect 3424 142128 3476 142180
rect 183744 142128 183796 142180
rect 120724 142060 120776 142112
rect 126060 142060 126112 142112
rect 157340 142060 157392 142112
rect 189448 142060 189500 142112
rect 117964 141924 118016 141976
rect 126796 141924 126848 141976
rect 184204 141924 184256 141976
rect 187240 141924 187292 141976
rect 183192 141856 183244 141908
rect 193772 141856 193824 141908
rect 115480 141788 115532 141840
rect 127348 141788 127400 141840
rect 181996 141788 182048 141840
rect 196348 141788 196400 141840
rect 114100 141720 114152 141772
rect 126244 141720 126296 141772
rect 179512 141720 179564 141772
rect 180340 141720 180392 141772
rect 197728 141720 197780 141772
rect 119896 141652 119948 141704
rect 138112 141652 138164 141704
rect 175188 141652 175240 141704
rect 193496 141652 193548 141704
rect 118148 141584 118200 141636
rect 146852 141584 146904 141636
rect 170772 141584 170824 141636
rect 192024 141584 192076 141636
rect 120816 141516 120868 141568
rect 152372 141516 152424 141568
rect 169116 141516 169168 141568
rect 192300 141516 192352 141568
rect 120908 141448 120960 141500
rect 153292 141448 153344 141500
rect 167460 141448 167512 141500
rect 192208 141448 192260 141500
rect 119436 141380 119488 141432
rect 153752 141380 153804 141432
rect 157156 141380 157208 141432
rect 189356 141380 189408 141432
rect 119804 141312 119856 141364
rect 123484 141312 123536 141364
rect 116860 141244 116912 141296
rect 125508 141244 125560 141296
rect 185032 141176 185084 141228
rect 185676 141176 185728 141228
rect 126060 141108 126112 141160
rect 129464 141108 129516 141160
rect 184756 141108 184808 141160
rect 190920 141108 190972 141160
rect 117964 141040 118016 141092
rect 179512 141040 179564 141092
rect 17224 140972 17276 141024
rect 185032 140972 185084 141024
rect 8944 140904 8996 140956
rect 182916 140904 182968 140956
rect 185860 140904 185912 140956
rect 191196 140904 191248 140956
rect 126796 140836 126848 140888
rect 129464 140836 129516 140888
rect 327724 140836 327776 140888
rect 464344 140768 464396 140820
rect 119528 140700 119580 140752
rect 119344 140632 119396 140684
rect 124772 140632 124824 140684
rect 128360 140700 128412 140752
rect 129280 140700 129332 140752
rect 131304 140700 131356 140752
rect 132316 140700 132368 140752
rect 129004 140632 129056 140684
rect 113640 140564 113692 140616
rect 129096 140564 129148 140616
rect 121000 140496 121052 140548
rect 146944 140700 146996 140752
rect 178040 140700 178092 140752
rect 178960 140700 179012 140752
rect 146760 140632 146812 140684
rect 173900 140632 173952 140684
rect 179144 140632 179196 140684
rect 119252 140428 119304 140480
rect 171140 140564 171192 140616
rect 190828 140700 190880 140752
rect 184480 140564 184532 140616
rect 193956 140564 194008 140616
rect 178132 140496 178184 140548
rect 178592 140496 178644 140548
rect 179972 140496 180024 140548
rect 193588 140496 193640 140548
rect 179052 140428 179104 140480
rect 196624 140428 196676 140480
rect 119436 140360 119488 140412
rect 148232 140360 148284 140412
rect 171232 140360 171284 140412
rect 189724 140360 189776 140412
rect 116400 140292 116452 140344
rect 145564 140292 145616 140344
rect 169852 140292 169904 140344
rect 189540 140292 189592 140344
rect 116584 140224 116636 140276
rect 147956 140224 148008 140276
rect 171324 140224 171376 140276
rect 192392 140224 192444 140276
rect 117872 140156 117924 140208
rect 149428 140156 149480 140208
rect 169944 140156 169996 140208
rect 185584 140156 185636 140208
rect 116768 140088 116820 140140
rect 150072 140088 150124 140140
rect 170864 140088 170916 140140
rect 192576 140156 192628 140208
rect 119160 140020 119212 140072
rect 126152 140020 126204 140072
rect 126612 140020 126664 140072
rect 184664 140020 184716 140072
rect 185676 140020 185728 140072
rect 196440 140020 196492 140072
rect 120632 139952 120684 140004
rect 129188 139952 129240 140004
rect 129464 139952 129516 140004
rect 183008 139952 183060 140004
rect 189908 139952 189960 140004
rect 124772 139884 124824 139936
rect 184572 139884 184624 139936
rect 189632 139884 189684 139936
rect 119804 139816 119856 139868
rect 126520 139816 126572 139868
rect 185584 139816 185636 139868
rect 192668 139816 192720 139868
rect 118056 139680 118108 139732
rect 124864 139680 124916 139732
rect 128820 139544 128872 139596
rect 178040 139544 178092 139596
rect 181628 139544 181680 139596
rect 188620 139544 188672 139596
rect 127532 139476 127584 139528
rect 181812 139476 181864 139528
rect 124864 139408 124916 139460
rect 181904 139408 181956 139460
rect 183284 139408 183336 139460
rect 189816 139408 189868 139460
rect 126152 139340 126204 139392
rect 126428 139340 126480 139392
rect 3516 137912 3568 137964
rect 117964 137912 118016 137964
rect 3148 111732 3200 111784
rect 31024 111732 31076 111784
rect 3516 97928 3568 97980
rect 120540 97928 120592 97980
rect 107292 89088 107344 89140
rect 107384 88884 107436 88936
rect 464344 86912 464396 86964
rect 580172 86912 580224 86964
rect 121920 81200 121972 81252
rect 122196 81200 122248 81252
rect 123116 81064 123168 81116
rect 121644 80996 121696 81048
rect 108304 80860 108356 80912
rect 120724 80860 120776 80912
rect 71780 80656 71832 80708
rect 108396 80656 108448 80708
rect 116584 80656 116636 80708
rect 120724 80656 120776 80708
rect 130016 80656 130068 80708
rect 131672 80656 131724 80708
rect 187424 81200 187476 81252
rect 187516 81064 187568 81116
rect 192668 81064 192720 81116
rect 131856 80656 131908 80708
rect 106740 80384 106792 80436
rect 107016 80384 107068 80436
rect 130752 80316 130804 80368
rect 107016 80248 107068 80300
rect 107200 80248 107252 80300
rect 131856 80248 131908 80300
rect 131764 80180 131816 80232
rect 131580 80112 131632 80164
rect 119160 80044 119212 80096
rect 130752 80044 130804 80096
rect 131672 80044 131724 80096
rect 130660 79976 130712 80028
rect 130476 79908 130528 79960
rect 132638 79908 132690 79960
rect 132822 79908 132874 79960
rect 133098 79908 133150 79960
rect 133282 79908 133334 79960
rect 133374 79908 133426 79960
rect 133466 79908 133518 79960
rect 133558 79908 133610 79960
rect 133742 79908 133794 79960
rect 133834 79908 133886 79960
rect 133926 79908 133978 79960
rect 134110 79908 134162 79960
rect 134386 79908 134438 79960
rect 134570 79908 134622 79960
rect 132132 79840 132184 79892
rect 132914 79840 132966 79892
rect 129464 79772 129516 79824
rect 133190 79840 133242 79892
rect 109868 79704 109920 79756
rect 131764 79704 131816 79756
rect 133144 79704 133196 79756
rect 116216 79636 116268 79688
rect 133512 79772 133564 79824
rect 133420 79704 133472 79756
rect 112352 79568 112404 79620
rect 122840 79568 122892 79620
rect 124128 79568 124180 79620
rect 113824 79500 113876 79552
rect 125600 79500 125652 79552
rect 106832 79432 106884 79484
rect 126244 79432 126296 79484
rect 133328 79636 133380 79688
rect 133052 79568 133104 79620
rect 133742 79772 133794 79824
rect 133788 79636 133840 79688
rect 132408 79500 132460 79552
rect 134018 79840 134070 79892
rect 134202 79840 134254 79892
rect 134294 79840 134346 79892
rect 134248 79704 134300 79756
rect 134156 79636 134208 79688
rect 134064 79568 134116 79620
rect 134432 79636 134484 79688
rect 134340 79568 134392 79620
rect 134754 79840 134806 79892
rect 134938 79908 134990 79960
rect 135214 79908 135266 79960
rect 135306 79908 135358 79960
rect 136134 79908 136186 79960
rect 136318 79908 136370 79960
rect 135950 79840 136002 79892
rect 135352 79772 135404 79824
rect 135674 79772 135726 79824
rect 135766 79772 135818 79824
rect 135168 79636 135220 79688
rect 135720 79636 135772 79688
rect 134708 79568 134760 79620
rect 135628 79568 135680 79620
rect 136226 79840 136278 79892
rect 136364 79772 136416 79824
rect 136272 79704 136324 79756
rect 135996 79636 136048 79688
rect 136180 79636 136232 79688
rect 134524 79500 134576 79552
rect 135076 79500 135128 79552
rect 135812 79500 135864 79552
rect 136686 79908 136738 79960
rect 136732 79704 136784 79756
rect 137146 79908 137198 79960
rect 137100 79704 137152 79756
rect 137422 79908 137474 79960
rect 137974 79908 138026 79960
rect 138066 79908 138118 79960
rect 138158 79908 138210 79960
rect 138250 79908 138302 79960
rect 137698 79840 137750 79892
rect 137284 79636 137336 79688
rect 137560 79636 137612 79688
rect 137882 79772 137934 79824
rect 138020 79772 138072 79824
rect 138112 79772 138164 79824
rect 138204 79704 138256 79756
rect 137836 79636 137888 79688
rect 136916 79568 136968 79620
rect 136456 79500 136508 79552
rect 138618 79908 138670 79960
rect 139262 79908 139314 79960
rect 139630 79908 139682 79960
rect 138802 79840 138854 79892
rect 139078 79840 139130 79892
rect 138572 79500 138624 79552
rect 139216 79636 139268 79688
rect 139308 79568 139360 79620
rect 139400 79568 139452 79620
rect 139860 79568 139912 79620
rect 139216 79500 139268 79552
rect 140044 79500 140096 79552
rect 140366 79908 140418 79960
rect 140458 79908 140510 79960
rect 140550 79908 140602 79960
rect 141470 79908 141522 79960
rect 141562 79908 141614 79960
rect 142298 79908 142350 79960
rect 142574 79908 142626 79960
rect 142758 79908 142810 79960
rect 143402 79908 143454 79960
rect 140412 79772 140464 79824
rect 140228 79568 140280 79620
rect 141010 79840 141062 79892
rect 141654 79840 141706 79892
rect 141838 79840 141890 79892
rect 141424 79568 141476 79620
rect 140688 79500 140740 79552
rect 140872 79500 140924 79552
rect 141240 79500 141292 79552
rect 142022 79840 142074 79892
rect 143034 79840 143086 79892
rect 142620 79704 142672 79756
rect 142804 79704 142856 79756
rect 143678 79908 143730 79960
rect 144138 79908 144190 79960
rect 144230 79908 144282 79960
rect 144966 79908 145018 79960
rect 145334 79908 145386 79960
rect 145794 79908 145846 79960
rect 145886 79908 145938 79960
rect 146070 79908 146122 79960
rect 146254 79908 146306 79960
rect 146530 79908 146582 79960
rect 143954 79840 144006 79892
rect 143862 79772 143914 79824
rect 141884 79636 141936 79688
rect 141976 79636 142028 79688
rect 142252 79636 142304 79688
rect 142160 79432 142212 79484
rect 142712 79568 142764 79620
rect 143080 79568 143132 79620
rect 143448 79704 143500 79756
rect 143540 79704 143592 79756
rect 143356 79636 143408 79688
rect 143908 79636 143960 79688
rect 144598 79840 144650 79892
rect 144874 79840 144926 79892
rect 144184 79772 144236 79824
rect 144322 79772 144374 79824
rect 144414 79772 144466 79824
rect 144506 79772 144558 79824
rect 144092 79568 144144 79620
rect 144276 79568 144328 79620
rect 143264 79500 143316 79552
rect 143816 79500 143868 79552
rect 143080 79432 143132 79484
rect 143724 79432 143776 79484
rect 144736 79636 144788 79688
rect 144828 79568 144880 79620
rect 145426 79840 145478 79892
rect 145702 79840 145754 79892
rect 145748 79704 145800 79756
rect 145840 79704 145892 79756
rect 145472 79636 145524 79688
rect 145656 79636 145708 79688
rect 146024 79636 146076 79688
rect 146116 79636 146168 79688
rect 146346 79840 146398 79892
rect 146438 79840 146490 79892
rect 146300 79704 146352 79756
rect 146392 79704 146444 79756
rect 146576 79704 146628 79756
rect 146806 79908 146858 79960
rect 146990 79908 147042 79960
rect 147082 79908 147134 79960
rect 147174 79908 147226 79960
rect 147358 79908 147410 79960
rect 147818 79908 147870 79960
rect 148002 79908 148054 79960
rect 148094 79908 148146 79960
rect 148186 79908 148238 79960
rect 148738 79908 148790 79960
rect 147036 79772 147088 79824
rect 147450 79840 147502 79892
rect 147220 79772 147272 79824
rect 147312 79772 147364 79824
rect 147404 79704 147456 79756
rect 146668 79636 146720 79688
rect 146852 79636 146904 79688
rect 144644 79500 144696 79552
rect 144552 79432 144604 79484
rect 147128 79432 147180 79484
rect 148048 79704 148100 79756
rect 148278 79840 148330 79892
rect 148370 79840 148422 79892
rect 148554 79840 148606 79892
rect 147956 79636 148008 79688
rect 148140 79636 148192 79688
rect 148324 79636 148376 79688
rect 149198 79908 149250 79960
rect 149842 79908 149894 79960
rect 150118 79908 150170 79960
rect 150302 79908 150354 79960
rect 148830 79840 148882 79892
rect 149290 79840 149342 79892
rect 149382 79840 149434 79892
rect 148692 79772 148744 79824
rect 148600 79704 148652 79756
rect 149244 79704 149296 79756
rect 147864 79568 147916 79620
rect 148692 79568 148744 79620
rect 148508 79500 148560 79552
rect 148876 79432 148928 79484
rect 111156 79364 111208 79416
rect 131764 79364 131816 79416
rect 131856 79364 131908 79416
rect 142988 79364 143040 79416
rect 150026 79840 150078 79892
rect 150256 79772 150308 79824
rect 150670 79908 150722 79960
rect 150946 79908 150998 79960
rect 151130 79840 151182 79892
rect 150348 79704 150400 79756
rect 150164 79636 150216 79688
rect 151406 79908 151458 79960
rect 151498 79840 151550 79892
rect 186780 80996 186832 81048
rect 200764 80928 200816 80980
rect 187424 80860 187476 80912
rect 206192 80860 206244 80912
rect 234620 80860 234672 80912
rect 186780 80792 186832 80844
rect 252560 80792 252612 80844
rect 178776 80588 178828 80640
rect 188160 80724 188212 80776
rect 270500 80724 270552 80776
rect 195152 80656 195204 80708
rect 358820 80656 358872 80708
rect 177764 80452 177816 80504
rect 179604 80384 179656 80436
rect 152050 79908 152102 79960
rect 153062 79908 153114 79960
rect 153154 79908 153206 79960
rect 153246 79908 153298 79960
rect 152694 79840 152746 79892
rect 151314 79772 151366 79824
rect 150532 79568 150584 79620
rect 150716 79568 150768 79620
rect 151452 79704 151504 79756
rect 151360 79636 151412 79688
rect 151268 79568 151320 79620
rect 152556 79568 152608 79620
rect 149980 79432 150032 79484
rect 149704 79364 149756 79416
rect 149888 79364 149940 79416
rect 150900 79500 150952 79552
rect 152280 79500 152332 79552
rect 150808 79432 150860 79484
rect 151544 79432 151596 79484
rect 151728 79432 151780 79484
rect 104900 79296 104952 79348
rect 106004 79296 106056 79348
rect 109776 79296 109828 79348
rect 132316 79296 132368 79348
rect 133236 79296 133288 79348
rect 135536 79296 135588 79348
rect 138296 79296 138348 79348
rect 138940 79296 138992 79348
rect 123668 79228 123720 79280
rect 149244 79296 149296 79348
rect 119344 79160 119396 79212
rect 141332 79160 141384 79212
rect 147956 79228 148008 79280
rect 151452 79228 151504 79280
rect 152096 79432 152148 79484
rect 152832 79432 152884 79484
rect 152648 79364 152700 79416
rect 152188 79296 152240 79348
rect 153108 79772 153160 79824
rect 153200 79704 153252 79756
rect 153430 79908 153482 79960
rect 178040 80316 178092 80368
rect 153706 79840 153758 79892
rect 154074 79840 154126 79892
rect 154166 79840 154218 79892
rect 154120 79704 154172 79756
rect 153936 79636 153988 79688
rect 154304 79636 154356 79688
rect 154534 79908 154586 79960
rect 154626 79908 154678 79960
rect 154718 79908 154770 79960
rect 154672 79704 154724 79756
rect 155178 79908 155230 79960
rect 155270 79908 155322 79960
rect 155730 79908 155782 79960
rect 155914 79908 155966 79960
rect 156098 79908 156150 79960
rect 156282 79908 156334 79960
rect 156466 79908 156518 79960
rect 156558 79908 156610 79960
rect 156834 79908 156886 79960
rect 156926 79908 156978 79960
rect 157294 79908 157346 79960
rect 157662 79908 157714 79960
rect 154488 79636 154540 79688
rect 155040 79636 155092 79688
rect 120632 79092 120684 79144
rect 142988 79160 143040 79212
rect 155270 79772 155322 79824
rect 155638 79772 155690 79824
rect 155224 79636 155276 79688
rect 155684 79568 155736 79620
rect 155316 79432 155368 79484
rect 156282 79772 156334 79824
rect 156512 79568 156564 79620
rect 156696 79568 156748 79620
rect 156328 79500 156380 79552
rect 156420 79432 156472 79484
rect 156052 79364 156104 79416
rect 156972 79772 157024 79824
rect 156972 79500 157024 79552
rect 157570 79772 157622 79824
rect 157616 79500 157668 79552
rect 158306 79908 158358 79960
rect 159042 79908 159094 79960
rect 159134 79908 159186 79960
rect 159594 79908 159646 79960
rect 160422 79908 160474 79960
rect 160514 79908 160566 79960
rect 160882 79908 160934 79960
rect 161066 79908 161118 79960
rect 161158 79908 161210 79960
rect 161250 79908 161302 79960
rect 158214 79840 158266 79892
rect 158030 79772 158082 79824
rect 158490 79840 158542 79892
rect 158076 79636 158128 79688
rect 158352 79636 158404 79688
rect 158674 79840 158726 79892
rect 158766 79840 158818 79892
rect 158536 79568 158588 79620
rect 158628 79568 158680 79620
rect 157524 79432 157576 79484
rect 157800 79432 157852 79484
rect 158904 79500 158956 79552
rect 159778 79840 159830 79892
rect 159548 79772 159600 79824
rect 160376 79772 160428 79824
rect 160468 79704 160520 79756
rect 160698 79840 160750 79892
rect 160790 79840 160842 79892
rect 160744 79704 160796 79756
rect 160836 79636 160888 79688
rect 160652 79568 160704 79620
rect 160928 79568 160980 79620
rect 161342 79772 161394 79824
rect 161112 79704 161164 79756
rect 161204 79636 161256 79688
rect 161296 79568 161348 79620
rect 161618 79908 161670 79960
rect 161986 79908 162038 79960
rect 162170 79908 162222 79960
rect 162998 79908 163050 79960
rect 163090 79908 163142 79960
rect 163366 79908 163418 79960
rect 163734 79908 163786 79960
rect 164010 79908 164062 79960
rect 164102 79908 164154 79960
rect 164470 79908 164522 79960
rect 164838 79908 164890 79960
rect 164930 79908 164982 79960
rect 165206 79908 165258 79960
rect 161664 79772 161716 79824
rect 161894 79772 161946 79824
rect 162354 79840 162406 79892
rect 162538 79840 162590 79892
rect 162630 79840 162682 79892
rect 162814 79840 162866 79892
rect 161848 79636 161900 79688
rect 162216 79636 162268 79688
rect 162584 79704 162636 79756
rect 162676 79704 162728 79756
rect 161940 79568 161992 79620
rect 162400 79568 162452 79620
rect 159640 79500 159692 79552
rect 159916 79500 159968 79552
rect 159088 79432 159140 79484
rect 159364 79432 159416 79484
rect 159732 79364 159784 79416
rect 161572 79364 161624 79416
rect 163274 79840 163326 79892
rect 162952 79704 163004 79756
rect 163182 79772 163234 79824
rect 163044 79568 163096 79620
rect 163228 79636 163280 79688
rect 163826 79840 163878 79892
rect 163458 79772 163510 79824
rect 163320 79568 163372 79620
rect 163136 79500 163188 79552
rect 163780 79568 163832 79620
rect 163872 79568 163924 79620
rect 164194 79840 164246 79892
rect 164286 79840 164338 79892
rect 164102 79772 164154 79824
rect 164332 79704 164384 79756
rect 164240 79568 164292 79620
rect 165482 79840 165534 79892
rect 165252 79772 165304 79824
rect 164930 79704 164982 79756
rect 164792 79636 164844 79688
rect 163596 79432 163648 79484
rect 164884 79568 164936 79620
rect 165068 79568 165120 79620
rect 165344 79568 165396 79620
rect 164424 79500 164476 79552
rect 164700 79500 164752 79552
rect 164976 79500 165028 79552
rect 165942 79908 165994 79960
rect 166126 79908 166178 79960
rect 166218 79908 166270 79960
rect 166310 79908 166362 79960
rect 166402 79908 166454 79960
rect 166494 79908 166546 79960
rect 165758 79772 165810 79824
rect 165804 79636 165856 79688
rect 166080 79772 166132 79824
rect 166172 79704 166224 79756
rect 166770 79840 166822 79892
rect 166862 79840 166914 79892
rect 166448 79704 166500 79756
rect 166632 79636 166684 79688
rect 166356 79568 166408 79620
rect 167000 79568 167052 79620
rect 165988 79500 166040 79552
rect 166724 79500 166776 79552
rect 165068 79432 165120 79484
rect 165620 79432 165672 79484
rect 167230 79908 167282 79960
rect 167690 79908 167742 79960
rect 167184 79568 167236 79620
rect 168334 79908 168386 79960
rect 168426 79908 168478 79960
rect 168518 79908 168570 79960
rect 168886 79908 168938 79960
rect 169070 79908 169122 79960
rect 168288 79772 168340 79824
rect 168426 79772 168478 79824
rect 168610 79772 168662 79824
rect 168564 79568 168616 79620
rect 168656 79568 168708 79620
rect 168978 79840 169030 79892
rect 169116 79772 169168 79824
rect 169714 79908 169766 79960
rect 169806 79908 169858 79960
rect 169990 79908 170042 79960
rect 169346 79840 169398 79892
rect 169622 79840 169674 79892
rect 169208 79568 169260 79620
rect 169392 79568 169444 79620
rect 168012 79500 168064 79552
rect 168840 79500 168892 79552
rect 169898 79840 169950 79892
rect 169852 79704 169904 79756
rect 169668 79568 169720 79620
rect 169760 79500 169812 79552
rect 169392 79432 169444 79484
rect 170036 79636 170088 79688
rect 170266 79908 170318 79960
rect 170358 79840 170410 79892
rect 170542 79908 170594 79960
rect 170726 79908 170778 79960
rect 171094 79908 171146 79960
rect 171186 79908 171238 79960
rect 170910 79840 170962 79892
rect 170220 79568 170272 79620
rect 170312 79500 170364 79552
rect 170404 79500 170456 79552
rect 170864 79636 170916 79688
rect 171370 79908 171422 79960
rect 171324 79772 171376 79824
rect 171232 79704 171284 79756
rect 179880 80248 179932 80300
rect 179328 80180 179380 80232
rect 171738 79908 171790 79960
rect 172014 79908 172066 79960
rect 172382 79908 172434 79960
rect 172842 79908 172894 79960
rect 172934 79908 172986 79960
rect 173026 79908 173078 79960
rect 173210 79908 173262 79960
rect 173302 79908 173354 79960
rect 173394 79908 173446 79960
rect 171048 79636 171100 79688
rect 171140 79568 171192 79620
rect 171416 79636 171468 79688
rect 172060 79772 172112 79824
rect 172336 79772 172388 79824
rect 172980 79772 173032 79824
rect 172796 79704 172848 79756
rect 173256 79772 173308 79824
rect 173348 79772 173400 79824
rect 173670 79908 173722 79960
rect 173762 79908 173814 79960
rect 173578 79840 173630 79892
rect 173716 79772 173768 79824
rect 178500 80112 178552 80164
rect 177764 80044 177816 80096
rect 181168 80044 181220 80096
rect 238760 80044 238812 80096
rect 173946 79908 173998 79960
rect 174406 79908 174458 79960
rect 174590 79908 174642 79960
rect 174682 79908 174734 79960
rect 174774 79908 174826 79960
rect 173624 79704 173676 79756
rect 173808 79704 173860 79756
rect 174222 79840 174274 79892
rect 174498 79840 174550 79892
rect 173900 79636 173952 79688
rect 174360 79772 174412 79824
rect 174958 79840 175010 79892
rect 175050 79840 175102 79892
rect 174728 79772 174780 79824
rect 174866 79772 174918 79824
rect 174636 79704 174688 79756
rect 175004 79704 175056 79756
rect 175510 79908 175562 79960
rect 175970 79908 176022 79960
rect 177856 79976 177908 80028
rect 175464 79772 175516 79824
rect 175602 79772 175654 79824
rect 175694 79772 175746 79824
rect 174544 79636 174596 79688
rect 174820 79636 174872 79688
rect 175096 79636 175148 79688
rect 175648 79636 175700 79688
rect 154764 79296 154816 79348
rect 164424 79296 164476 79348
rect 171692 79364 171744 79416
rect 174176 79432 174228 79484
rect 175280 79568 175332 79620
rect 176154 79840 176206 79892
rect 176246 79840 176298 79892
rect 177074 79908 177126 79960
rect 175924 79636 175976 79688
rect 176430 79772 176482 79824
rect 176200 79704 176252 79756
rect 176292 79704 176344 79756
rect 176384 79636 176436 79688
rect 176798 79840 176850 79892
rect 177856 79840 177908 79892
rect 176706 79772 176758 79824
rect 177580 79772 177632 79824
rect 178592 79976 178644 80028
rect 178224 79704 178276 79756
rect 191288 79704 191340 79756
rect 176108 79568 176160 79620
rect 178132 79636 178184 79688
rect 189816 79636 189868 79688
rect 177488 79568 177540 79620
rect 190736 79568 190788 79620
rect 175372 79500 175424 79552
rect 175832 79500 175884 79552
rect 176752 79500 176804 79552
rect 178776 79500 178828 79552
rect 178040 79432 178092 79484
rect 194048 79432 194100 79484
rect 163964 79228 164016 79280
rect 165712 79228 165764 79280
rect 165896 79228 165948 79280
rect 174360 79296 174412 79348
rect 177764 79296 177816 79348
rect 306380 79364 306432 79416
rect 189908 79296 189960 79348
rect 167368 79160 167420 79212
rect 193864 79228 193916 79280
rect 196808 79160 196860 79212
rect 119252 79024 119304 79076
rect 147404 79092 147456 79144
rect 160652 79092 160704 79144
rect 118056 78956 118108 79008
rect 147220 79024 147272 79076
rect 157616 79024 157668 79076
rect 173164 79024 173216 79076
rect 192944 79092 192996 79144
rect 173808 79024 173860 79076
rect 192024 79024 192076 79076
rect 324320 79296 324372 79348
rect 142160 78956 142212 79008
rect 147864 78956 147916 79008
rect 168104 78956 168156 79008
rect 168288 78956 168340 79008
rect 201868 78956 201920 79008
rect 117596 78888 117648 78940
rect 140504 78888 140556 78940
rect 141332 78888 141384 78940
rect 145380 78888 145432 78940
rect 148692 78888 148744 78940
rect 117872 78820 117924 78872
rect 157616 78888 157668 78940
rect 157800 78888 157852 78940
rect 163964 78888 164016 78940
rect 169024 78888 169076 78940
rect 169208 78888 169260 78940
rect 170864 78888 170916 78940
rect 171508 78888 171560 78940
rect 172152 78888 172204 78940
rect 172612 78888 172664 78940
rect 181076 78888 181128 78940
rect 288440 78888 288492 78940
rect 130108 78752 130160 78804
rect 140044 78752 140096 78804
rect 180892 78820 180944 78872
rect 186320 78820 186372 78872
rect 186964 78820 187016 78872
rect 480260 78820 480312 78872
rect 149060 78752 149112 78804
rect 150072 78752 150124 78804
rect 152004 78752 152056 78804
rect 152188 78752 152240 78804
rect 170312 78752 170364 78804
rect 172612 78752 172664 78804
rect 173164 78752 173216 78804
rect 173808 78752 173860 78804
rect 173992 78752 174044 78804
rect 178224 78752 178276 78804
rect 186412 78752 186464 78804
rect 187056 78752 187108 78804
rect 483020 78752 483072 78804
rect 131856 78684 131908 78736
rect 137560 78684 137612 78736
rect 140964 78684 141016 78736
rect 141332 78684 141384 78736
rect 146852 78684 146904 78736
rect 179512 78684 179564 78736
rect 187700 78684 187752 78736
rect 188344 78684 188396 78736
rect 500960 78684 501012 78736
rect 120080 78616 120132 78668
rect 121368 78616 121420 78668
rect 132040 78616 132092 78668
rect 133696 78616 133748 78668
rect 133880 78616 133932 78668
rect 138388 78616 138440 78668
rect 138572 78616 138624 78668
rect 138848 78616 138900 78668
rect 139124 78616 139176 78668
rect 140504 78616 140556 78668
rect 146300 78616 146352 78668
rect 148968 78616 149020 78668
rect 152004 78616 152056 78668
rect 152372 78616 152424 78668
rect 153292 78616 153344 78668
rect 154120 78616 154172 78668
rect 165804 78616 165856 78668
rect 196256 78616 196308 78668
rect 196624 78616 196676 78668
rect 102140 78548 102192 78600
rect 102784 78548 102836 78600
rect 134064 78548 134116 78600
rect 137560 78548 137612 78600
rect 143356 78548 143408 78600
rect 147220 78548 147272 78600
rect 150532 78548 150584 78600
rect 164424 78548 164476 78600
rect 130844 78480 130896 78532
rect 133880 78480 133932 78532
rect 104072 78412 104124 78464
rect 130476 78412 130528 78464
rect 132592 78344 132644 78396
rect 142620 78480 142672 78532
rect 142988 78480 143040 78532
rect 169668 78548 169720 78600
rect 170312 78480 170364 78532
rect 171876 78480 171928 78532
rect 172244 78480 172296 78532
rect 181444 78548 181496 78600
rect 192852 78548 192904 78600
rect 186320 78480 186372 78532
rect 137100 78412 137152 78464
rect 142068 78412 142120 78464
rect 153752 78412 153804 78464
rect 154488 78412 154540 78464
rect 158812 78412 158864 78464
rect 163412 78412 163464 78464
rect 170036 78412 170088 78464
rect 186412 78412 186464 78464
rect 139124 78344 139176 78396
rect 139308 78344 139360 78396
rect 140964 78344 141016 78396
rect 141424 78344 141476 78396
rect 142620 78344 142672 78396
rect 142988 78344 143040 78396
rect 143540 78344 143592 78396
rect 163228 78344 163280 78396
rect 164148 78344 164200 78396
rect 165896 78344 165948 78396
rect 166172 78344 166224 78396
rect 167000 78344 167052 78396
rect 183100 78344 183152 78396
rect 205824 78344 205876 78396
rect 206192 78344 206244 78396
rect 57980 78276 58032 78328
rect 107292 78276 107344 78328
rect 122196 78276 122248 78328
rect 148508 78276 148560 78328
rect 167460 78276 167512 78328
rect 253204 78276 253256 78328
rect 46940 78208 46992 78260
rect 107200 78208 107252 78260
rect 123392 78208 123444 78260
rect 20720 78140 20772 78192
rect 102140 78140 102192 78192
rect 6920 78072 6972 78124
rect 107108 78072 107160 78124
rect 107384 78072 107436 78124
rect 2780 78004 2832 78056
rect 104072 78004 104124 78056
rect 2872 77936 2924 77988
rect 108580 77936 108632 77988
rect 130200 78140 130252 78192
rect 133880 78140 133932 78192
rect 137560 78140 137612 78192
rect 138296 78208 138348 78260
rect 144092 78208 144144 78260
rect 150624 78208 150676 78260
rect 151176 78208 151228 78260
rect 160928 78208 160980 78260
rect 166172 78208 166224 78260
rect 169852 78208 169904 78260
rect 170864 78208 170916 78260
rect 337384 78208 337436 78260
rect 148324 78140 148376 78192
rect 152556 78140 152608 78192
rect 153016 78140 153068 78192
rect 161480 78140 161532 78192
rect 162032 78140 162084 78192
rect 400864 78140 400916 78192
rect 123024 78072 123076 78124
rect 143448 78072 143500 78124
rect 149704 78072 149756 78124
rect 183652 78072 183704 78124
rect 196256 78072 196308 78124
rect 429200 78072 429252 78124
rect 113640 78004 113692 78056
rect 129832 78004 129884 78056
rect 131856 78004 131908 78056
rect 132500 77936 132552 77988
rect 137100 77936 137152 77988
rect 153200 77936 153252 77988
rect 153660 77936 153712 77988
rect 156420 77936 156472 77988
rect 161480 77936 161532 77988
rect 131028 77868 131080 77920
rect 142528 77868 142580 77920
rect 148416 77868 148468 77920
rect 148784 77868 148836 77920
rect 107384 77800 107436 77852
rect 129464 77800 129516 77852
rect 129556 77800 129608 77852
rect 134432 77800 134484 77852
rect 131948 77732 132000 77784
rect 150440 77800 150492 77852
rect 151452 77800 151504 77852
rect 157432 77800 157484 77852
rect 157800 77800 157852 77852
rect 159364 77732 159416 77784
rect 173992 78004 174044 78056
rect 174176 78004 174228 78056
rect 178960 78004 179012 78056
rect 180800 78004 180852 78056
rect 415492 78004 415544 78056
rect 169484 77936 169536 77988
rect 169760 77936 169812 77988
rect 177396 77936 177448 77988
rect 177856 77936 177908 77988
rect 162952 77868 163004 77920
rect 177212 77868 177264 77920
rect 163504 77800 163556 77852
rect 178776 77800 178828 77852
rect 165252 77732 165304 77784
rect 422300 77936 422352 77988
rect 181536 77868 181588 77920
rect 194140 77868 194192 77920
rect 107292 77664 107344 77716
rect 136824 77664 136876 77716
rect 137100 77664 137152 77716
rect 142344 77664 142396 77716
rect 169852 77664 169904 77716
rect 171140 77664 171192 77716
rect 187516 77664 187568 77716
rect 131212 77596 131264 77648
rect 132316 77596 132368 77648
rect 139860 77596 139912 77648
rect 156144 77596 156196 77648
rect 162216 77596 162268 77648
rect 131764 77528 131816 77580
rect 142252 77528 142304 77580
rect 164608 77528 164660 77580
rect 180800 77528 180852 77580
rect 107200 77460 107252 77512
rect 136088 77460 136140 77512
rect 137008 77460 137060 77512
rect 137376 77460 137428 77512
rect 164056 77460 164108 77512
rect 178868 77460 178920 77512
rect 134064 77392 134116 77444
rect 137560 77392 137612 77444
rect 138112 77392 138164 77444
rect 146024 77392 146076 77444
rect 158352 77392 158404 77444
rect 163504 77392 163556 77444
rect 164700 77392 164752 77444
rect 165068 77392 165120 77444
rect 181444 77392 181496 77444
rect 130200 77324 130252 77376
rect 133604 77324 133656 77376
rect 154856 77324 154908 77376
rect 158628 77324 158680 77376
rect 160744 77324 160796 77376
rect 161388 77324 161440 77376
rect 161664 77324 161716 77376
rect 167644 77324 167696 77376
rect 169944 77324 169996 77376
rect 170680 77324 170732 77376
rect 176384 77324 176436 77376
rect 177304 77324 177356 77376
rect 179328 77324 179380 77376
rect 132776 77256 132828 77308
rect 105544 77188 105596 77240
rect 105820 77188 105872 77240
rect 124864 77188 124916 77240
rect 125600 77188 125652 77240
rect 133144 77188 133196 77240
rect 162216 77256 162268 77308
rect 177488 77256 177540 77308
rect 137468 77188 137520 77240
rect 159456 77188 159508 77240
rect 161664 77188 161716 77240
rect 172796 77188 172848 77240
rect 205824 77188 205876 77240
rect 206100 77188 206152 77240
rect 122380 77120 122432 77172
rect 144460 77120 144512 77172
rect 145656 77120 145708 77172
rect 156696 77120 156748 77172
rect 156880 77120 156932 77172
rect 161020 77120 161072 77172
rect 191196 77120 191248 77172
rect 191748 77120 191800 77172
rect 118976 77052 119028 77104
rect 108488 76984 108540 77036
rect 106004 76916 106056 76968
rect 130292 76916 130344 76968
rect 118516 76848 118568 76900
rect 130384 76848 130436 76900
rect 72424 76712 72476 76764
rect 106924 76780 106976 76832
rect 132684 76916 132736 76968
rect 133144 76984 133196 77036
rect 141884 76984 141936 77036
rect 147772 77052 147824 77104
rect 147956 77052 148008 77104
rect 159824 77052 159876 77104
rect 189632 77052 189684 77104
rect 152648 76984 152700 77036
rect 133328 76916 133380 76968
rect 144184 76916 144236 76968
rect 151820 76916 151872 76968
rect 133604 76848 133656 76900
rect 134064 76780 134116 76832
rect 136916 76780 136968 76832
rect 149428 76848 149480 76900
rect 149980 76848 150032 76900
rect 148784 76780 148836 76832
rect 119436 76712 119488 76764
rect 148600 76712 148652 76764
rect 177948 76984 178000 77036
rect 205916 76984 205968 77036
rect 155500 76916 155552 76968
rect 179328 76916 179380 76968
rect 170220 76848 170272 76900
rect 170588 76848 170640 76900
rect 192576 76848 192628 76900
rect 170680 76780 170732 76832
rect 192760 76780 192812 76832
rect 260840 76712 260892 76764
rect 64144 76644 64196 76696
rect 106004 76644 106056 76696
rect 117412 76644 117464 76696
rect 132776 76644 132828 76696
rect 134524 76644 134576 76696
rect 139032 76644 139084 76696
rect 143540 76644 143592 76696
rect 144092 76644 144144 76696
rect 148324 76644 148376 76696
rect 148692 76644 148744 76696
rect 149336 76644 149388 76696
rect 52460 76576 52512 76628
rect 135812 76576 135864 76628
rect 149612 76576 149664 76628
rect 150256 76576 150308 76628
rect 161756 76644 161808 76696
rect 161940 76644 161992 76696
rect 162860 76644 162912 76696
rect 163044 76644 163096 76696
rect 167184 76644 167236 76696
rect 169116 76644 169168 76696
rect 170864 76644 170916 76696
rect 189540 76644 189592 76696
rect 189632 76644 189684 76696
rect 353300 76644 353352 76696
rect 181444 76576 181496 76628
rect 191748 76576 191800 76628
rect 367100 76576 367152 76628
rect 35900 76508 35952 76560
rect 135260 76508 135312 76560
rect 151268 76508 151320 76560
rect 203708 76508 203760 76560
rect 205824 76508 205876 76560
rect 509884 76508 509936 76560
rect 126244 76440 126296 76492
rect 133144 76440 133196 76492
rect 133328 76440 133380 76492
rect 140412 76440 140464 76492
rect 161756 76440 161808 76492
rect 162400 76440 162452 76492
rect 162860 76440 162912 76492
rect 164240 76440 164292 76492
rect 168564 76440 168616 76492
rect 168748 76440 168800 76492
rect 169024 76440 169076 76492
rect 178684 76440 178736 76492
rect 112444 76372 112496 76424
rect 146668 76372 146720 76424
rect 153936 76372 153988 76424
rect 160836 76372 160888 76424
rect 161296 76372 161348 76424
rect 168840 76372 168892 76424
rect 169208 76372 169260 76424
rect 105544 76304 105596 76356
rect 132776 76304 132828 76356
rect 141056 76304 141108 76356
rect 171968 76304 172020 76356
rect 189724 76304 189776 76356
rect 140136 76236 140188 76288
rect 133144 76168 133196 76220
rect 141700 76168 141752 76220
rect 164240 76168 164292 76220
rect 165804 76168 165856 76220
rect 164608 76032 164660 76084
rect 164884 76032 164936 76084
rect 172704 76032 172756 76084
rect 173624 76032 173676 76084
rect 158628 75964 158680 76016
rect 180064 75964 180116 76016
rect 289820 75964 289872 76016
rect 104900 75828 104952 75880
rect 110788 75828 110840 75880
rect 111064 75828 111116 75880
rect 146024 75896 146076 75948
rect 146944 75896 146996 75948
rect 164516 75896 164568 75948
rect 165160 75896 165212 75948
rect 167092 75896 167144 75948
rect 167736 75896 167788 75948
rect 171968 75896 172020 75948
rect 172152 75896 172204 75948
rect 179328 75896 179380 75948
rect 296720 75896 296772 75948
rect 139400 75828 139452 75880
rect 144460 75828 144512 75880
rect 151084 75828 151136 75880
rect 163596 75828 163648 75880
rect 163872 75828 163924 75880
rect 198464 75828 198516 75880
rect 107016 75760 107068 75812
rect 138020 75760 138072 75812
rect 164424 75760 164476 75812
rect 165436 75760 165488 75812
rect 165804 75760 165856 75812
rect 166080 75760 166132 75812
rect 166908 75760 166960 75812
rect 167184 75760 167236 75812
rect 171416 75760 171468 75812
rect 171968 75760 172020 75812
rect 115388 75692 115440 75744
rect 146392 75692 146444 75744
rect 154304 75692 154356 75744
rect 163136 75692 163188 75744
rect 166264 75692 166316 75744
rect 170404 75692 170456 75744
rect 171048 75692 171100 75744
rect 187976 75760 188028 75812
rect 178500 75692 178552 75744
rect 183560 75692 183612 75744
rect 111064 75624 111116 75676
rect 139952 75624 140004 75676
rect 146760 75624 146812 75676
rect 182824 75624 182876 75676
rect 108672 75556 108724 75608
rect 135444 75556 135496 75608
rect 153936 75556 153988 75608
rect 187700 75556 187752 75608
rect 115204 75488 115256 75540
rect 117412 75488 117464 75540
rect 121276 75488 121328 75540
rect 146576 75488 146628 75540
rect 147956 75488 148008 75540
rect 148048 75488 148100 75540
rect 201500 75488 201552 75540
rect 122564 75420 122616 75472
rect 145196 75420 145248 75472
rect 150348 75420 150400 75472
rect 216680 75420 216732 75472
rect 81440 75352 81492 75404
rect 138664 75352 138716 75404
rect 166356 75352 166408 75404
rect 166908 75352 166960 75404
rect 172980 75352 173032 75404
rect 480904 75352 480956 75404
rect 67640 75284 67692 75336
rect 137652 75284 137704 75336
rect 145104 75284 145156 75336
rect 145748 75284 145800 75336
rect 172244 75284 172296 75336
rect 506480 75284 506532 75336
rect 22744 75216 22796 75268
rect 132408 75216 132460 75268
rect 135812 75216 135864 75268
rect 136364 75216 136416 75268
rect 139492 75216 139544 75268
rect 140320 75216 140372 75268
rect 153200 75216 153252 75268
rect 153844 75216 153896 75268
rect 158904 75216 158956 75268
rect 159180 75216 159232 75268
rect 172336 75216 172388 75268
rect 511264 75216 511316 75268
rect 7564 75148 7616 75200
rect 120080 75148 120132 75200
rect 122288 75148 122340 75200
rect 145564 75148 145616 75200
rect 168012 75148 168064 75200
rect 130016 75080 130068 75132
rect 131028 75080 131080 75132
rect 162676 75080 162728 75132
rect 164792 75080 164844 75132
rect 168748 75080 168800 75132
rect 169300 75080 169352 75132
rect 178040 75148 178092 75200
rect 549260 75148 549312 75200
rect 154120 75012 154172 75064
rect 154396 75012 154448 75064
rect 176844 75080 176896 75132
rect 177120 75080 177172 75132
rect 177764 75080 177816 75132
rect 180064 75012 180116 75064
rect 205732 75012 205784 75064
rect 154304 74944 154356 74996
rect 180800 74944 180852 74996
rect 135444 74876 135496 74928
rect 136548 74876 136600 74928
rect 177028 74876 177080 74928
rect 177488 74876 177540 74928
rect 132960 74740 133012 74792
rect 133512 74740 133564 74792
rect 109960 74468 110012 74520
rect 144000 74536 144052 74588
rect 175832 74536 175884 74588
rect 176108 74536 176160 74588
rect 142252 74468 142304 74520
rect 143172 74468 143224 74520
rect 153292 74468 153344 74520
rect 154028 74468 154080 74520
rect 166908 74468 166960 74520
rect 200948 74468 201000 74520
rect 110052 74400 110104 74452
rect 144644 74400 144696 74452
rect 153384 74400 153436 74452
rect 188620 74400 188672 74452
rect 269120 74400 269172 74452
rect 112904 74332 112956 74384
rect 111524 74264 111576 74316
rect 141516 74264 141568 74316
rect 143172 74332 143224 74384
rect 143448 74332 143500 74384
rect 171508 74332 171560 74384
rect 172152 74332 172204 74384
rect 172888 74332 172940 74384
rect 173532 74332 173584 74384
rect 198280 74332 198332 74384
rect 144920 74264 144972 74316
rect 172520 74264 172572 74316
rect 173440 74264 173492 74316
rect 196992 74264 197044 74316
rect 111432 74196 111484 74248
rect 143908 74196 143960 74248
rect 147128 74196 147180 74248
rect 150992 74196 151044 74248
rect 237380 74196 237432 74248
rect 100208 74128 100260 74180
rect 133788 74128 133840 74180
rect 141516 74128 141568 74180
rect 144552 74128 144604 74180
rect 152372 74128 152424 74180
rect 255320 74128 255372 74180
rect 104164 74060 104216 74112
rect 135536 74060 135588 74112
rect 153476 74060 153528 74112
rect 284300 74060 284352 74112
rect 93860 73992 93912 74044
rect 104900 73992 104952 74044
rect 123208 73992 123260 74044
rect 153292 73992 153344 74044
rect 155592 73992 155644 74044
rect 297364 73992 297416 74044
rect 104256 73924 104308 73976
rect 134156 73924 134208 73976
rect 134616 73924 134668 73976
rect 161664 73924 161716 73976
rect 347780 73924 347832 73976
rect 54484 73856 54536 73908
rect 107568 73856 107620 73908
rect 112812 73856 112864 73908
rect 142252 73856 142304 73908
rect 152740 73856 152792 73908
rect 261484 73856 261536 73908
rect 269764 73856 269816 73908
rect 465172 73856 465224 73908
rect 21364 73788 21416 73840
rect 100208 73788 100260 73840
rect 112996 73788 113048 73840
rect 142528 73788 142580 73840
rect 151728 73788 151780 73840
rect 248420 73788 248472 73840
rect 253204 73788 253256 73840
rect 449900 73788 449952 73840
rect 114192 73720 114244 73772
rect 142988 73720 143040 73772
rect 155040 73720 155092 73772
rect 155684 73720 155736 73772
rect 172520 73720 172572 73772
rect 173348 73720 173400 73772
rect 107568 73652 107620 73704
rect 136456 73652 136508 73704
rect 172152 73652 172204 73704
rect 192392 73720 192444 73772
rect 104256 73312 104308 73364
rect 104624 73312 104676 73364
rect 111340 73176 111392 73228
rect 114560 73176 114612 73228
rect 115848 73176 115900 73228
rect 110236 73108 110288 73160
rect 144092 73108 144144 73160
rect 157340 73108 157392 73160
rect 158260 73108 158312 73160
rect 160376 73108 160428 73160
rect 161112 73108 161164 73160
rect 167828 73108 167880 73160
rect 168012 73108 168064 73160
rect 202328 73108 202380 73160
rect 327724 73108 327776 73160
rect 580172 73108 580224 73160
rect 123760 73040 123812 73092
rect 149336 73040 149388 73092
rect 149888 73040 149940 73092
rect 157524 73040 157576 73092
rect 158536 73040 158588 73092
rect 165988 73040 166040 73092
rect 198096 73040 198148 73092
rect 206284 73040 206336 73092
rect 119988 72972 120040 73024
rect 152004 72972 152056 73024
rect 155684 72972 155736 73024
rect 190092 72972 190144 73024
rect 106096 72904 106148 72956
rect 139124 72904 139176 72956
rect 144000 72904 144052 72956
rect 144276 72904 144328 72956
rect 163412 72904 163464 72956
rect 163688 72904 163740 72956
rect 164700 72904 164752 72956
rect 165436 72904 165488 72956
rect 199476 72904 199528 72956
rect 107476 72836 107528 72888
rect 138572 72836 138624 72888
rect 155960 72836 156012 72888
rect 156972 72836 157024 72888
rect 167000 72836 167052 72888
rect 202420 72836 202472 72888
rect 111616 72768 111668 72820
rect 143080 72768 143132 72820
rect 156604 72768 156656 72820
rect 311164 72768 311216 72820
rect 104440 72700 104492 72752
rect 130660 72700 130712 72752
rect 157248 72700 157300 72752
rect 318800 72700 318852 72752
rect 115848 72632 115900 72684
rect 141148 72632 141200 72684
rect 157708 72632 157760 72684
rect 324964 72632 325016 72684
rect 70400 72564 70452 72616
rect 137836 72564 137888 72616
rect 157616 72564 157668 72616
rect 332600 72564 332652 72616
rect 23480 72496 23532 72548
rect 100300 72496 100352 72548
rect 14464 72428 14516 72480
rect 104440 72428 104492 72480
rect 123944 72496 123996 72548
rect 149520 72496 149572 72548
rect 149888 72496 149940 72548
rect 166172 72496 166224 72548
rect 368480 72496 368532 72548
rect 116492 72428 116544 72480
rect 141608 72428 141660 72480
rect 158260 72428 158312 72480
rect 191104 72428 191156 72480
rect 202420 72428 202472 72480
rect 446404 72428 446456 72480
rect 122748 72360 122800 72412
rect 129924 72360 129976 72412
rect 132500 72360 132552 72412
rect 145012 72360 145064 72412
rect 145380 72360 145432 72412
rect 158536 72360 158588 72412
rect 190000 72360 190052 72412
rect 167000 72292 167052 72344
rect 168104 72292 168156 72344
rect 176108 72292 176160 72344
rect 204536 72292 204588 72344
rect 134340 72224 134392 72276
rect 152004 72224 152056 72276
rect 152832 72224 152884 72276
rect 161112 72224 161164 72276
rect 187240 72224 187292 72276
rect 134340 72088 134392 72140
rect 135168 72088 135220 72140
rect 175924 72088 175976 72140
rect 176292 72088 176344 72140
rect 128912 71952 128964 72004
rect 133236 71952 133288 72004
rect 115940 71748 115992 71800
rect 116492 71748 116544 71800
rect 124956 71748 125008 71800
rect 126244 71748 126296 71800
rect 127348 71748 127400 71800
rect 122104 71680 122156 71732
rect 122840 71680 122892 71732
rect 123300 71680 123352 71732
rect 127440 71680 127492 71732
rect 3516 71612 3568 71664
rect 8944 71612 8996 71664
rect 99380 71612 99432 71664
rect 100392 71612 100444 71664
rect 151912 71680 151964 71732
rect 156420 71680 156472 71732
rect 156696 71680 156748 71732
rect 159640 71680 159692 71732
rect 160008 71680 160060 71732
rect 160836 71680 160888 71732
rect 161296 71680 161348 71732
rect 161940 71680 161992 71732
rect 162584 71680 162636 71732
rect 183652 71680 183704 71732
rect 204444 71680 204496 71732
rect 134432 71612 134484 71664
rect 141424 71612 141476 71664
rect 143080 71612 143132 71664
rect 151360 71612 151412 71664
rect 151544 71612 151596 71664
rect 117504 71544 117556 71596
rect 127348 71544 127400 71596
rect 127808 71544 127860 71596
rect 158812 71612 158864 71664
rect 159732 71612 159784 71664
rect 160284 71612 160336 71664
rect 161020 71612 161072 71664
rect 194968 71612 195020 71664
rect 162584 71544 162636 71596
rect 196440 71544 196492 71596
rect 116952 71476 117004 71528
rect 149796 71476 149848 71528
rect 158812 71476 158864 71528
rect 159364 71476 159416 71528
rect 169668 71476 169720 71528
rect 203524 71476 203576 71528
rect 108764 71408 108816 71460
rect 140596 71408 140648 71460
rect 162124 71408 162176 71460
rect 196900 71408 196952 71460
rect 120816 71340 120868 71392
rect 152464 71340 152516 71392
rect 161296 71340 161348 71392
rect 194232 71340 194284 71392
rect 119068 71272 119120 71324
rect 121000 71204 121052 71256
rect 162400 71272 162452 71324
rect 195428 71272 195480 71324
rect 27620 71136 27672 71188
rect 99380 71136 99432 71188
rect 108948 71136 109000 71188
rect 138204 71136 138256 71188
rect 139216 71136 139268 71188
rect 151268 71204 151320 71256
rect 159732 71204 159784 71256
rect 192300 71204 192352 71256
rect 151360 71136 151412 71188
rect 151912 71136 151964 71188
rect 152648 71136 152700 71188
rect 166632 71136 166684 71188
rect 166816 71136 166868 71188
rect 187148 71136 187200 71188
rect 26240 71068 26292 71120
rect 102140 71068 102192 71120
rect 113456 71068 113508 71120
rect 140412 71068 140464 71120
rect 148968 71068 149020 71120
rect 179420 71068 179472 71120
rect 179512 71068 179564 71120
rect 185032 71068 185084 71120
rect 45560 71000 45612 71052
rect 135996 71000 136048 71052
rect 160468 71000 160520 71052
rect 188344 71068 188396 71120
rect 196624 71068 196676 71120
rect 204444 71068 204496 71120
rect 218060 71068 218112 71120
rect 354680 71000 354732 71052
rect 117688 70932 117740 70984
rect 136824 70932 136876 70984
rect 142896 70932 142948 70984
rect 160008 70932 160060 70984
rect 114284 70864 114336 70916
rect 128360 70864 128412 70916
rect 137100 70864 137152 70916
rect 160100 70864 160152 70916
rect 160744 70864 160796 70916
rect 180892 70932 180944 70984
rect 188344 70932 188396 70984
rect 193956 70864 194008 70916
rect 102140 70796 102192 70848
rect 103060 70796 103112 70848
rect 129556 70796 129608 70848
rect 144276 70796 144328 70848
rect 147128 70796 147180 70848
rect 189172 70728 189224 70780
rect 189356 70728 189408 70780
rect 142528 70660 142580 70712
rect 142988 70660 143040 70712
rect 107660 70388 107712 70440
rect 108764 70388 108816 70440
rect 119620 70320 119672 70372
rect 153200 70320 153252 70372
rect 153844 70320 153896 70372
rect 167184 70320 167236 70372
rect 168104 70320 168156 70372
rect 202144 70320 202196 70372
rect 121736 70252 121788 70304
rect 155224 70252 155276 70304
rect 167276 70252 167328 70304
rect 167828 70252 167880 70304
rect 202236 70252 202288 70304
rect 120448 70184 120500 70236
rect 153660 70184 153712 70236
rect 154212 70184 154264 70236
rect 162492 70184 162544 70236
rect 196532 70184 196584 70236
rect 120908 70116 120960 70168
rect 154120 70116 154172 70168
rect 164976 70116 165028 70168
rect 199568 70116 199620 70168
rect 122012 70048 122064 70100
rect 46204 69708 46256 69760
rect 102968 69708 103020 69760
rect 131580 69980 131632 70032
rect 144552 70048 144604 70100
rect 146300 70048 146352 70100
rect 165344 70048 165396 70100
rect 199660 70048 199712 70100
rect 153568 69980 153620 70032
rect 153936 69980 153988 70032
rect 163872 69980 163924 70032
rect 113548 69912 113600 69964
rect 142528 69912 142580 69964
rect 143264 69912 143316 69964
rect 164332 69912 164384 69964
rect 164976 69912 165028 69964
rect 165160 69980 165212 70032
rect 199384 69980 199436 70032
rect 198188 69912 198240 69964
rect 112720 69844 112772 69896
rect 139492 69844 139544 69896
rect 161664 69844 161716 69896
rect 162492 69844 162544 69896
rect 164516 69844 164568 69896
rect 165344 69844 165396 69896
rect 165896 69844 165948 69896
rect 166632 69844 166684 69896
rect 200856 69844 200908 69896
rect 115020 69776 115072 69828
rect 142160 69776 142212 69828
rect 142620 69776 142672 69828
rect 163044 69776 163096 69828
rect 163872 69776 163924 69828
rect 164608 69776 164660 69828
rect 165160 69776 165212 69828
rect 169116 69776 169168 69828
rect 201776 69776 201828 69828
rect 202788 69776 202840 69828
rect 115572 69708 115624 69760
rect 138112 69708 138164 69760
rect 138572 69708 138624 69760
rect 139492 69708 139544 69760
rect 140320 69708 140372 69760
rect 164424 69708 164476 69760
rect 188528 69708 188580 69760
rect 423772 69708 423824 69760
rect 18604 69640 18656 69692
rect 119804 69640 119856 69692
rect 128452 69640 128504 69692
rect 142436 69640 142488 69692
rect 147956 69640 148008 69692
rect 181536 69640 181588 69692
rect 202788 69640 202840 69692
rect 448520 69640 448572 69692
rect 103152 69572 103204 69624
rect 130200 69572 130252 69624
rect 103520 69504 103572 69556
rect 108488 69504 108540 69556
rect 109040 68960 109092 69012
rect 110972 68960 111024 69012
rect 118332 68960 118384 69012
rect 152280 68960 152332 69012
rect 152556 68960 152608 69012
rect 167092 68960 167144 69012
rect 168288 68960 168340 69012
rect 202052 68960 202104 69012
rect 117228 68892 117280 68944
rect 151176 68892 151228 68944
rect 161480 68892 161532 68944
rect 189172 68892 189224 68944
rect 108856 68824 108908 68876
rect 142344 68824 142396 68876
rect 142712 68824 142764 68876
rect 176936 68824 176988 68876
rect 199384 68824 199436 68876
rect 104624 68756 104676 68808
rect 136088 68756 136140 68808
rect 163596 68756 163648 68808
rect 183008 68756 183060 68808
rect 183468 68756 183520 68808
rect 89720 68552 89772 68604
rect 105728 68552 105780 68604
rect 131028 68552 131080 68604
rect 135260 68552 135312 68604
rect 85580 68484 85632 68536
rect 106096 68484 106148 68536
rect 120080 68484 120132 68536
rect 141792 68484 141844 68536
rect 78680 68416 78732 68468
rect 107476 68416 107528 68468
rect 118608 68416 118660 68468
rect 141240 68416 141292 68468
rect 149888 68416 149940 68468
rect 220820 68416 220872 68468
rect 75920 68348 75972 68400
rect 107016 68348 107068 68400
rect 117320 68348 117372 68400
rect 140964 68348 141016 68400
rect 189172 68348 189224 68400
rect 302240 68348 302292 68400
rect 48320 68280 48372 68332
rect 104624 68280 104676 68332
rect 113180 68280 113232 68332
rect 140780 68280 140832 68332
rect 186688 68280 186740 68332
rect 504364 68280 504416 68332
rect 183468 67668 183520 67720
rect 332692 67668 332744 67720
rect 199384 67600 199436 67652
rect 560944 67600 560996 67652
rect 104348 67532 104400 67584
rect 138480 67532 138532 67584
rect 144920 67532 144972 67584
rect 147220 67532 147272 67584
rect 165804 67532 165856 67584
rect 200396 67532 200448 67584
rect 201408 67532 201460 67584
rect 114008 67464 114060 67516
rect 139860 67464 139912 67516
rect 110144 67396 110196 67448
rect 118608 67396 118660 67448
rect 92480 67124 92532 67176
rect 105636 67124 105688 67176
rect 93952 67056 94004 67108
rect 112536 67056 112588 67108
rect 80060 66988 80112 67040
rect 104348 66988 104400 67040
rect 106280 66988 106332 67040
rect 139584 66988 139636 67040
rect 102140 66920 102192 66972
rect 139676 66920 139728 66972
rect 164792 66920 164844 66972
rect 389180 66920 389232 66972
rect 99380 66852 99432 66904
rect 139768 66852 139820 66904
rect 201408 66852 201460 66904
rect 432604 66852 432656 66904
rect 140780 66240 140832 66292
rect 142160 66240 142212 66292
rect 189172 66240 189224 66292
rect 539600 66240 539652 66292
rect 102232 66172 102284 66224
rect 103244 66172 103296 66224
rect 134340 66172 134392 66224
rect 144000 66172 144052 66224
rect 148416 66172 148468 66224
rect 159088 66172 159140 66224
rect 190920 66172 190972 66224
rect 191748 66172 191800 66224
rect 98000 65560 98052 65612
rect 111064 65560 111116 65612
rect 148784 65560 148836 65612
rect 207020 65560 207072 65612
rect 35992 65492 36044 65544
rect 102232 65492 102284 65544
rect 146484 65492 146536 65544
rect 183560 65492 183612 65544
rect 191748 65492 191800 65544
rect 346400 65492 346452 65544
rect 139400 64880 139452 64932
rect 142160 64880 142212 64932
rect 102232 64812 102284 64864
rect 103336 64812 103388 64864
rect 137192 64812 137244 64864
rect 168840 64812 168892 64864
rect 203064 64812 203116 64864
rect 149704 64268 149756 64320
rect 224960 64268 225012 64320
rect 62120 64200 62172 64252
rect 102232 64200 102284 64252
rect 152832 64200 152884 64252
rect 256700 64200 256752 64252
rect 4160 64132 4212 64184
rect 132500 64132 132552 64184
rect 150532 64132 150584 64184
rect 183008 64132 183060 64184
rect 203064 64132 203116 64184
rect 472624 64132 472676 64184
rect 104716 63452 104768 63504
rect 132776 63452 132828 63504
rect 158996 63452 159048 63504
rect 193220 63452 193272 63504
rect 88340 62840 88392 62892
rect 138388 62840 138440 62892
rect 193220 62840 193272 62892
rect 340880 62840 340932 62892
rect 10324 62772 10376 62824
rect 104716 62772 104768 62824
rect 160192 62772 160244 62824
rect 357440 62772 357492 62824
rect 102232 62024 102284 62076
rect 103428 62024 103480 62076
rect 135812 62024 135864 62076
rect 162952 62024 163004 62076
rect 197360 62024 197412 62076
rect 197544 62024 197596 62076
rect 166356 61956 166408 62008
rect 197636 61956 197688 62008
rect 135352 61888 135404 61940
rect 142988 61888 143040 61940
rect 176844 61888 176896 61940
rect 196072 61888 196124 61940
rect 172704 61820 172756 61872
rect 186964 61820 187016 61872
rect 144644 61480 144696 61532
rect 149704 61480 149756 61532
rect 52552 61412 52604 61464
rect 102232 61412 102284 61464
rect 197360 61412 197412 61464
rect 394700 61412 394752 61464
rect 42800 61344 42852 61396
rect 135720 61344 135772 61396
rect 197636 61344 197688 61396
rect 198372 61344 198424 61396
rect 396080 61344 396132 61396
rect 186964 60800 187016 60852
rect 529940 60800 529992 60852
rect 196072 60732 196124 60784
rect 574744 60732 574796 60784
rect 99472 60664 99524 60716
rect 100576 60664 100628 60716
rect 133604 60664 133656 60716
rect 158904 60664 158956 60716
rect 193312 60664 193364 60716
rect 194508 60664 194560 60716
rect 104808 60596 104860 60648
rect 137468 60596 137520 60648
rect 149796 60188 149848 60240
rect 223580 60188 223632 60240
rect 145196 60120 145248 60172
rect 147312 60120 147364 60172
rect 150808 60120 150860 60172
rect 245660 60120 245712 60172
rect 69020 60052 69072 60104
rect 104808 60052 104860 60104
rect 155316 60052 155368 60104
rect 299480 60052 299532 60104
rect 17960 59984 18012 60036
rect 99472 59984 99524 60036
rect 153108 59984 153160 60036
rect 186320 59984 186372 60036
rect 194508 59984 194560 60036
rect 345020 59984 345072 60036
rect 110420 59304 110472 59356
rect 115204 59304 115256 59356
rect 111800 59236 111852 59288
rect 112260 59236 112312 59288
rect 135996 59304 136048 59356
rect 147404 58692 147456 58744
rect 193312 58692 193364 58744
rect 49700 58624 49752 58676
rect 111800 58624 111852 58676
rect 170496 58624 170548 58676
rect 490012 58624 490064 58676
rect 168748 57876 168800 57928
rect 203432 57876 203484 57928
rect 204168 57876 204220 57928
rect 151452 57264 151504 57316
rect 233240 57264 233292 57316
rect 204168 57196 204220 57248
rect 473452 57196 473504 57248
rect 99472 56516 99524 56568
rect 100668 56516 100720 56568
rect 133420 56516 133472 56568
rect 63500 55904 63552 55956
rect 137008 55904 137060 55956
rect 147864 55904 147916 55956
rect 197360 55904 197412 55956
rect 12440 55836 12492 55888
rect 99472 55836 99524 55888
rect 148692 55836 148744 55888
rect 204260 55836 204312 55888
rect 138664 55224 138716 55276
rect 142344 55224 142396 55276
rect 168656 55156 168708 55208
rect 201684 55156 201736 55208
rect 202788 55156 202840 55208
rect 148140 54544 148192 54596
rect 209872 54544 209924 54596
rect 171048 54476 171100 54528
rect 486424 54476 486476 54528
rect 202788 53796 202840 53848
rect 464344 53796 464396 53848
rect 100484 53728 100536 53780
rect 133052 53728 133104 53780
rect 168564 53728 168616 53780
rect 203800 53728 203852 53780
rect 149244 53184 149296 53236
rect 215300 53184 215352 53236
rect 157984 53116 158036 53168
rect 333980 53116 334032 53168
rect 9680 53048 9732 53100
rect 100484 53048 100536 53100
rect 102232 53048 102284 53100
rect 113824 53048 113876 53100
rect 203800 53048 203852 53100
rect 466460 53048 466512 53100
rect 169208 52368 169260 52420
rect 202972 52368 203024 52420
rect 204168 52368 204220 52420
rect 145104 51824 145156 51876
rect 169024 51824 169076 51876
rect 155960 51756 156012 51808
rect 320180 51756 320232 51808
rect 147588 51688 147640 51740
rect 191840 51688 191892 51740
rect 204168 51688 204220 51740
rect 468484 51688 468536 51740
rect 100760 51008 100812 51060
rect 105544 51008 105596 51060
rect 176752 51008 176804 51060
rect 203064 51008 203116 51060
rect 204168 51008 204220 51060
rect 150164 50464 150216 50516
rect 218152 50464 218204 50516
rect 152740 50396 152792 50448
rect 259460 50396 259512 50448
rect 176660 50328 176712 50380
rect 578240 50328 578292 50380
rect 204168 49716 204220 49768
rect 569960 49716 570012 49768
rect 150256 49104 150308 49156
rect 222200 49104 222252 49156
rect 155224 49036 155276 49088
rect 285680 49036 285732 49088
rect 175280 48968 175332 49020
rect 556160 48968 556212 49020
rect 147772 47744 147824 47796
rect 201592 47744 201644 47796
rect 148600 47676 148652 47728
rect 208400 47676 208452 47728
rect 170588 47608 170640 47660
rect 488540 47608 488592 47660
rect 145012 47540 145064 47592
rect 168564 47540 168616 47592
rect 177672 47540 177724 47592
rect 582380 47540 582432 47592
rect 143816 46860 143868 46912
rect 147772 46860 147824 46912
rect 177488 46860 177540 46912
rect 204352 46860 204404 46912
rect 204720 46860 204772 46912
rect 151360 46384 151412 46436
rect 236000 46384 236052 46436
rect 154304 46316 154356 46368
rect 275284 46316 275336 46368
rect 168380 46248 168432 46300
rect 474740 46248 474792 46300
rect 204720 46180 204772 46232
rect 571984 46180 572036 46232
rect 161572 44956 161624 45008
rect 390560 44956 390612 45008
rect 172520 44888 172572 44940
rect 527180 44888 527232 44940
rect 60832 44820 60884 44872
rect 137928 44820 137980 44872
rect 174636 44820 174688 44872
rect 542360 44820 542412 44872
rect 156328 43528 156380 43580
rect 315304 43528 315356 43580
rect 163780 43460 163832 43512
rect 404360 43460 404412 43512
rect 162860 43392 162912 43444
rect 408500 43392 408552 43444
rect 138020 42576 138072 42628
rect 142252 42576 142304 42628
rect 155408 42304 155460 42356
rect 292672 42304 292724 42356
rect 164240 42236 164292 42288
rect 426440 42236 426492 42288
rect 166540 42168 166592 42220
rect 440332 42168 440384 42220
rect 171324 42100 171376 42152
rect 498292 42100 498344 42152
rect 77392 42032 77444 42084
rect 138848 42032 138900 42084
rect 173624 42032 173676 42084
rect 528560 42032 528612 42084
rect 148508 40944 148560 40996
rect 205640 40944 205692 40996
rect 157064 40876 157116 40928
rect 317420 40876 317472 40928
rect 165712 40808 165764 40860
rect 444380 40808 444432 40860
rect 173440 40740 173492 40792
rect 516140 40740 516192 40792
rect 13820 40672 13872 40724
rect 132868 40672 132920 40724
rect 176200 40672 176252 40724
rect 564532 40672 564584 40724
rect 152648 39584 152700 39636
rect 251180 39584 251232 39636
rect 160744 39516 160796 39568
rect 361580 39516 361632 39568
rect 168472 39448 168524 39500
rect 463700 39448 463752 39500
rect 167000 39380 167052 39432
rect 462320 39380 462372 39432
rect 31760 39312 31812 39364
rect 134248 39312 134300 39364
rect 173532 39312 173584 39364
rect 520280 39312 520332 39364
rect 154672 38156 154724 38208
rect 293960 38156 294012 38208
rect 158812 38088 158864 38140
rect 351920 38088 351972 38140
rect 167828 38020 167880 38072
rect 448612 38020 448664 38072
rect 170680 37952 170732 38004
rect 481640 37952 481692 38004
rect 38660 37884 38712 37936
rect 135628 37884 135680 37936
rect 143724 37884 143776 37936
rect 154580 37884 154632 37936
rect 174728 37884 174780 37936
rect 538220 37884 538272 37936
rect 149060 36728 149112 36780
rect 226340 36728 226392 36780
rect 155500 36660 155552 36712
rect 299572 36660 299624 36712
rect 170772 36592 170824 36644
rect 484400 36592 484452 36644
rect 176108 36524 176160 36576
rect 552020 36524 552072 36576
rect 156880 35436 156932 35488
rect 310520 35436 310572 35488
rect 159732 35368 159784 35420
rect 342260 35368 342312 35420
rect 167920 35300 167972 35352
rect 454040 35300 454092 35352
rect 171784 35232 171836 35284
rect 502340 35232 502392 35284
rect 53840 35164 53892 35216
rect 135444 35164 135496 35216
rect 144920 35164 144972 35216
rect 167000 35164 167052 35216
rect 177764 35164 177816 35216
rect 571340 35164 571392 35216
rect 152556 34008 152608 34060
rect 251272 34008 251324 34060
rect 163872 33940 163924 33992
rect 391940 33940 391992 33992
rect 165068 33872 165120 33924
rect 410524 33872 410576 33924
rect 170864 33804 170916 33856
rect 491300 33804 491352 33856
rect 177856 33736 177908 33788
rect 576860 33736 576912 33788
rect 178960 33056 179012 33108
rect 580172 33056 580224 33108
rect 154212 32580 154264 32632
rect 267832 32580 267884 32632
rect 161020 32512 161072 32564
rect 357532 32512 357584 32564
rect 166724 32444 166776 32496
rect 431960 32444 432012 32496
rect 174820 32376 174872 32428
rect 539692 32376 539744 32428
rect 148876 31356 148928 31408
rect 198740 31356 198792 31408
rect 157156 31288 157208 31340
rect 303620 31288 303672 31340
rect 163688 31220 163740 31272
rect 340972 31220 341024 31272
rect 164976 31152 165028 31204
rect 409880 31152 409932 31204
rect 183100 31084 183152 31136
rect 443000 31084 443052 31136
rect 44272 31016 44324 31068
rect 135536 31016 135588 31068
rect 169852 31016 169904 31068
rect 495440 31016 495492 31068
rect 158260 29860 158312 29912
rect 321560 29860 321612 29912
rect 167736 29792 167788 29844
rect 375380 29792 375432 29844
rect 166632 29724 166684 29776
rect 434720 29724 434772 29776
rect 177304 29656 177356 29708
rect 554780 29656 554832 29708
rect 175372 29588 175424 29640
rect 558184 29588 558236 29640
rect 143632 28908 143684 28960
rect 144920 28908 144972 28960
rect 151268 28500 151320 28552
rect 242992 28500 243044 28552
rect 159824 28432 159876 28484
rect 339500 28432 339552 28484
rect 162032 28364 162084 28416
rect 379520 28364 379572 28416
rect 168012 28296 168064 28348
rect 456892 28296 456944 28348
rect 171968 28228 172020 28280
rect 506572 28228 506624 28280
rect 162308 27072 162360 27124
rect 374092 27072 374144 27124
rect 178868 27004 178920 27056
rect 407120 27004 407172 27056
rect 172152 26936 172204 26988
rect 509240 26936 509292 26988
rect 173716 26868 173768 26920
rect 524420 26868 524472 26920
rect 154028 25780 154080 25832
rect 278780 25780 278832 25832
rect 162400 25712 162452 25764
rect 382372 25712 382424 25764
rect 165252 25644 165304 25696
rect 425060 25644 425112 25696
rect 172244 25576 172296 25628
rect 513380 25576 513432 25628
rect 173256 25508 173308 25560
rect 531412 25508 531464 25560
rect 154120 24284 154172 24336
rect 282920 24284 282972 24336
rect 163964 24216 164016 24268
rect 398932 24216 398984 24268
rect 173164 24148 173216 24200
rect 522304 24148 522356 24200
rect 146208 24080 146260 24132
rect 173256 24080 173308 24132
rect 175004 24080 175056 24132
rect 546500 24080 546552 24132
rect 149980 22992 150032 23044
rect 219440 22992 219492 23044
rect 159916 22924 159968 22976
rect 350540 22924 350592 22976
rect 165160 22856 165212 22908
rect 416780 22856 416832 22908
rect 168196 22788 168248 22840
rect 460940 22788 460992 22840
rect 174912 22720 174964 22772
rect 534080 22720 534132 22772
rect 157800 21564 157852 21616
rect 322940 21564 322992 21616
rect 158352 21496 158404 21548
rect 329840 21496 329892 21548
rect 158444 21428 158496 21480
rect 336740 21428 336792 21480
rect 337384 21428 337436 21480
rect 471980 21428 472032 21480
rect 158720 21360 158772 21412
rect 343640 21360 343692 21412
rect 289084 20612 289136 20664
rect 579988 20612 580040 20664
rect 154396 20204 154448 20256
rect 273260 20204 273312 20256
rect 153752 20136 153804 20188
rect 280160 20136 280212 20188
rect 155776 20068 155828 20120
rect 291200 20068 291252 20120
rect 161204 20000 161256 20052
rect 372620 20000 372672 20052
rect 155684 19932 155736 19984
rect 287060 19932 287112 19984
rect 287704 19932 287756 19984
rect 518900 19932 518952 19984
rect 155868 18776 155920 18828
rect 300860 18776 300912 18828
rect 176292 18708 176344 18760
rect 522396 18708 522448 18760
rect 176384 18640 176436 18692
rect 567200 18640 567252 18692
rect 177948 18572 178000 18624
rect 574100 18572 574152 18624
rect 150624 17484 150676 17536
rect 241520 17484 241572 17536
rect 165528 17416 165580 17468
rect 418160 17416 418212 17468
rect 166816 17348 166868 17400
rect 441620 17348 441672 17400
rect 168104 17280 168156 17332
rect 445760 17280 445812 17332
rect 145564 17212 145616 17264
rect 164884 17212 164936 17264
rect 169668 17212 169720 17264
rect 477500 17212 477552 17264
rect 153016 16124 153068 16176
rect 259552 16124 259604 16176
rect 161112 16056 161164 16108
rect 361120 16056 361172 16108
rect 160100 15988 160152 16040
rect 364616 15988 364668 16040
rect 164148 15920 164200 15972
rect 397736 15920 397788 15972
rect 400864 15920 400916 15972
rect 478880 15920 478932 15972
rect 165344 15852 165396 15904
rect 420920 15852 420972 15904
rect 153936 14696 153988 14748
rect 272432 14696 272484 14748
rect 156788 14628 156840 14680
rect 314660 14628 314712 14680
rect 179328 14560 179380 14612
rect 394240 14560 394292 14612
rect 164056 14492 164108 14544
rect 407212 14492 407264 14544
rect 171876 14424 171928 14476
rect 503720 14424 503772 14476
rect 153844 13336 153896 13388
rect 276020 13336 276072 13388
rect 158536 13268 158588 13320
rect 324412 13268 324464 13320
rect 178776 13200 178828 13252
rect 400864 13200 400916 13252
rect 165436 13132 165488 13184
rect 414296 13132 414348 13184
rect 172060 13064 172112 13116
rect 511264 13064 511316 13116
rect 150900 11908 150952 11960
rect 245200 11908 245252 11960
rect 162676 11840 162728 11892
rect 386696 11840 386748 11892
rect 165620 11772 165672 11824
rect 439136 11772 439188 11824
rect 175096 11704 175148 11756
rect 548616 11704 548668 11756
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 152464 10548 152516 10600
rect 258264 10548 258316 10600
rect 156696 10480 156748 10532
rect 307944 10480 307996 10532
rect 162492 10412 162544 10464
rect 385960 10412 386012 10464
rect 162768 10344 162820 10396
rect 390652 10344 390704 10396
rect 87512 10276 87564 10328
rect 138112 10276 138164 10328
rect 170956 10276 171008 10328
rect 493048 10276 493100 10328
rect 151176 9256 151228 9308
rect 234712 9256 234764 9308
rect 158628 9188 158680 9240
rect 329196 9188 329248 9240
rect 161388 9120 161440 9172
rect 365812 9120 365864 9172
rect 166908 9052 166960 9104
rect 432052 9052 432104 9104
rect 176476 8984 176528 9036
rect 556160 8984 556212 9036
rect 105728 8916 105780 8968
rect 139860 8916 139912 8968
rect 143540 8916 143592 8968
rect 151912 8916 151964 8968
rect 185584 8916 185636 8968
rect 581000 8916 581052 8968
rect 149152 7760 149204 7812
rect 227536 7760 227588 7812
rect 160008 7692 160060 7744
rect 350448 7692 350500 7744
rect 168288 7624 168340 7676
rect 453396 7624 453448 7676
rect 30104 7556 30156 7608
rect 134156 7556 134208 7608
rect 175188 7556 175240 7608
rect 545488 7556 545540 7608
rect 3424 6808 3476 6860
rect 17224 6808 17276 6860
rect 576124 6808 576176 6860
rect 580172 6808 580224 6860
rect 156420 6400 156472 6452
rect 316224 6400 316276 6452
rect 161296 6332 161348 6384
rect 371700 6332 371752 6384
rect 169760 6264 169812 6316
rect 482836 6264 482888 6316
rect 176568 6196 176620 6248
rect 558552 6196 558604 6248
rect 175832 6128 175884 6180
rect 563244 6128 563296 6180
rect 152096 4972 152148 5024
rect 266544 4972 266596 5024
rect 162584 4904 162636 4956
rect 378876 4904 378928 4956
rect 170404 4836 170456 4888
rect 486332 4836 486384 4888
rect 173900 4768 173952 4820
rect 541992 4768 542044 4820
rect 142804 4156 142856 4208
rect 143540 4156 143592 4208
rect 572 4088 624 4140
rect 7564 4088 7616 4140
rect 15936 4088 15988 4140
rect 17316 4088 17368 4140
rect 73804 4088 73856 4140
rect 75184 4088 75236 4140
rect 127624 4088 127676 4140
rect 134524 4088 134576 4140
rect 146944 4088 146996 4140
rect 147404 4088 147456 4140
rect 169024 4088 169076 4140
rect 173164 4088 173216 4140
rect 196624 4088 196676 4140
rect 200304 4088 200356 4140
rect 301596 4088 301648 4140
rect 309048 4088 309100 4140
rect 315304 4088 315356 4140
rect 317328 4088 317380 4140
rect 324964 4088 325016 4140
rect 326804 4088 326856 4140
rect 382924 4088 382976 4140
rect 384764 4088 384816 4140
rect 450544 4088 450596 4140
rect 452108 4088 452160 4140
rect 489184 4088 489236 4140
rect 491116 4088 491168 4140
rect 1676 4020 1728 4072
rect 8944 4020 8996 4072
rect 147312 4020 147364 4072
rect 150716 4020 150768 4072
rect 151820 4020 151872 4072
rect 153016 4020 153068 4072
rect 130844 3952 130896 4004
rect 144736 3952 144788 4004
rect 149704 3952 149756 4004
rect 157800 3952 157852 4004
rect 45928 3884 45980 3936
rect 46204 3884 46256 3936
rect 124680 3884 124732 3936
rect 140872 3884 140924 3936
rect 149796 3884 149848 3936
rect 156604 3884 156656 3936
rect 156696 3884 156748 3936
rect 170772 3884 170824 3936
rect 112812 3816 112864 3868
rect 117412 3816 117464 3868
rect 125876 3816 125928 3868
rect 129924 3816 129976 3868
rect 130752 3816 130804 3868
rect 162492 3816 162544 3868
rect 91560 3748 91612 3800
rect 139492 3748 139544 3800
rect 147220 3748 147272 3800
rect 163688 3748 163740 3800
rect 85672 3680 85724 3732
rect 127624 3680 127676 3732
rect 66720 3612 66772 3664
rect 72424 3612 72476 3664
rect 83280 3612 83332 3664
rect 127716 3612 127768 3664
rect 19432 3544 19484 3596
rect 21364 3544 21416 3596
rect 44180 3544 44232 3596
rect 45100 3544 45152 3596
rect 51356 3544 51408 3596
rect 54484 3544 54536 3596
rect 59636 3544 59688 3596
rect 64144 3544 64196 3596
rect 69112 3544 69164 3596
rect 129832 3680 129884 3732
rect 127900 3612 127952 3664
rect 138204 3680 138256 3732
rect 147128 3680 147180 3732
rect 150624 3680 150676 3732
rect 150716 3680 150768 3732
rect 164516 3680 164568 3732
rect 137652 3612 137704 3664
rect 138664 3612 138716 3664
rect 147036 3612 147088 3664
rect 149520 3612 149572 3664
rect 151084 3612 151136 3664
rect 128176 3544 128228 3596
rect 130384 3544 130436 3596
rect 130936 3544 130988 3596
rect 166080 3680 166132 3732
rect 184204 3748 184256 3800
rect 210976 3748 211028 3800
rect 211804 3748 211856 3800
rect 181444 3680 181496 3732
rect 212172 3680 212224 3732
rect 234620 3748 234672 3800
rect 235816 3748 235868 3800
rect 247592 3680 247644 3732
rect 423772 3680 423824 3732
rect 424968 3680 425020 3732
rect 171968 3612 172020 3664
rect 189816 3612 189868 3664
rect 193220 3612 193272 3664
rect 203708 3612 203760 3664
rect 240508 3612 240560 3664
rect 247684 3612 247736 3664
rect 254676 3612 254728 3664
rect 261484 3612 261536 3664
rect 262956 3612 263008 3664
rect 299572 3612 299624 3664
rect 300768 3612 300820 3664
rect 311164 3612 311216 3664
rect 312636 3612 312688 3664
rect 164884 3544 164936 3596
rect 168380 3544 168432 3596
rect 173256 3544 173308 3596
rect 177856 3544 177908 3596
rect 180064 3544 180116 3596
rect 181536 3544 181588 3596
rect 182548 3544 182600 3596
rect 183008 3544 183060 3596
rect 190828 3544 190880 3596
rect 193864 3544 193916 3596
rect 196808 3544 196860 3596
rect 206284 3544 206336 3596
rect 403624 3544 403676 3596
rect 407120 3544 407172 3596
rect 408408 3544 408460 3596
rect 410524 3544 410576 3596
rect 411904 3544 411956 3596
rect 418804 3544 418856 3596
rect 420184 3544 420236 3596
rect 422944 3544 422996 3596
rect 423772 3544 423824 3596
rect 431960 3544 432012 3596
rect 433248 3544 433300 3596
rect 440240 3544 440292 3596
rect 441528 3544 441580 3596
rect 446404 3544 446456 3596
rect 447416 3544 447468 3596
rect 448612 3544 448664 3596
rect 449808 3544 449860 3596
rect 453304 3544 453356 3596
rect 497096 3544 497148 3596
rect 574744 3544 574796 3596
rect 576308 3544 576360 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 6460 3476 6512 3528
rect 8760 3408 8812 3460
rect 10324 3408 10376 3460
rect 17040 3408 17092 3460
rect 18604 3408 18656 3460
rect 27620 3408 27672 3460
rect 28540 3408 28592 3460
rect 33600 3408 33652 3460
rect 45928 3408 45980 3460
rect 52460 3408 52512 3460
rect 53380 3408 53432 3460
rect 56048 3408 56100 3460
rect 57244 3408 57296 3460
rect 60740 3408 60792 3460
rect 61660 3408 61712 3460
rect 65524 3408 65576 3460
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 123484 3476 123536 3528
rect 124956 3476 125008 3528
rect 126980 3476 127032 3528
rect 128452 3476 128504 3528
rect 131764 3340 131816 3392
rect 137284 3408 137336 3460
rect 148324 3408 148376 3460
rect 175464 3476 175516 3528
rect 458088 3476 458140 3528
rect 468484 3476 468536 3528
rect 469864 3476 469916 3528
rect 472624 3476 472676 3528
rect 473452 3476 473504 3528
rect 486424 3476 486476 3528
rect 487620 3476 487672 3528
rect 504364 3476 504416 3528
rect 505376 3476 505428 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 509884 3476 509936 3528
rect 518348 3476 518400 3528
rect 527916 3476 527968 3528
rect 533712 3476 533764 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 545764 3476 545816 3528
rect 551468 3476 551520 3528
rect 558184 3476 558236 3528
rect 559748 3476 559800 3528
rect 563704 3476 563756 3528
rect 565636 3476 565688 3528
rect 567844 3476 567896 3528
rect 569132 3476 569184 3528
rect 571984 3476 572036 3528
rect 573916 3476 573968 3528
rect 147404 3340 147456 3392
rect 176660 3408 176712 3460
rect 178684 3408 178736 3460
rect 468668 3408 468720 3460
rect 480904 3408 480956 3460
rect 521844 3408 521896 3460
rect 522396 3408 522448 3460
rect 560852 3408 560904 3460
rect 560944 3408 560996 3460
rect 572720 3408 572772 3460
rect 275284 3340 275336 3392
rect 277124 3340 277176 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 340880 3340 340932 3392
rect 342168 3340 342220 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 364984 3340 365036 3392
rect 367008 3340 367060 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 414664 3340 414716 3392
rect 416688 3340 416740 3392
rect 38384 3136 38436 3188
rect 39304 3136 39356 3188
rect 148416 3136 148468 3188
rect 154212 3136 154264 3188
rect 171784 3136 171836 3188
rect 174268 3136 174320 3188
rect 200764 3136 200816 3188
rect 203892 3136 203944 3188
rect 297364 3136 297416 3188
rect 298468 3136 298520 3188
rect 511356 3136 511408 3188
rect 514760 3136 514812 3188
rect 122288 3068 122340 3120
rect 124864 3068 124916 3120
rect 134156 3068 134208 3120
rect 136824 3068 136876 3120
rect 182824 3068 182876 3120
rect 184940 3068 184992 3120
rect 522304 3068 522356 3120
rect 524236 3068 524288 3120
rect 20628 3000 20680 3052
rect 22744 3000 22796 3052
rect 23020 3000 23072 3052
rect 25504 3000 25556 3052
rect 132960 3000 133012 3052
rect 141424 3000 141476 3052
rect 182916 3000 182968 3052
rect 189724 3000 189776 3052
rect 464344 3000 464396 3052
rect 466276 3000 466328 3052
rect 514024 3000 514076 3052
rect 515956 3000 516008 3052
rect 12348 2932 12400 2984
rect 14464 2932 14516 2984
rect 432604 2932 432656 2984
rect 434444 2932 434496 2984
rect 118792 2864 118844 2916
rect 122104 2864 122156 2916
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700534 8156 703520
rect 24320 700602 24348 703520
rect 24308 700596 24360 700602
rect 24308 700538 24360 700544
rect 8116 700528 8168 700534
rect 8116 700470 8168 700476
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683262 3464 684247
rect 3424 683256 3476 683262
rect 3424 683198 3476 683204
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 7564 514820 7616 514826
rect 3424 514762 3476 514768
rect 7564 514762 7616 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 2778 371376 2834 371385
rect 2778 371311 2780 371320
rect 2832 371311 2834 371320
rect 2780 371282 2832 371288
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3344 318850 3372 319223
rect 3332 318844 3384 318850
rect 3332 318786 3384 318792
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3436 265674 3464 475623
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 4804 371340 4856 371346
rect 4804 371282 4856 371288
rect 3514 358456 3570 358465
rect 3514 358391 3516 358400
rect 3568 358391 3570 358400
rect 3516 358362 3568 358368
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 305046 3556 306167
rect 3516 305040 3568 305046
rect 3516 304982 3568 304988
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 4816 268462 4844 371282
rect 7576 271250 7604 514762
rect 8944 358420 8996 358426
rect 8944 358362 8996 358368
rect 8956 273970 8984 358362
rect 40052 279478 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 279472 40092 279478
rect 40040 279414 40092 279420
rect 8944 273964 8996 273970
rect 8944 273906 8996 273912
rect 7564 271244 7616 271250
rect 7564 271186 7616 271192
rect 71792 269890 71820 702986
rect 89180 700738 89208 703520
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 105464 699718 105492 703520
rect 137848 700874 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700868 137888 700874
rect 137836 700810 137888 700816
rect 152464 700392 152516 700398
rect 152464 700334 152516 700340
rect 148324 700324 148376 700330
rect 148324 700266 148376 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 71780 269884 71832 269890
rect 71780 269826 71832 269832
rect 4804 268456 4856 268462
rect 4804 268398 4856 268404
rect 3424 265668 3476 265674
rect 3424 265610 3476 265616
rect 106936 264246 106964 699654
rect 146300 696992 146352 696998
rect 146300 696934 146352 696940
rect 143632 616888 143684 616894
rect 143632 616830 143684 616836
rect 142436 590708 142488 590714
rect 142436 590650 142488 590656
rect 139584 484424 139636 484430
rect 139584 484366 139636 484372
rect 138664 430636 138716 430642
rect 138664 430578 138716 430584
rect 135260 351960 135312 351966
rect 135260 351902 135312 351908
rect 134524 324352 134576 324358
rect 134524 324294 134576 324300
rect 133144 271924 133196 271930
rect 133144 271866 133196 271872
rect 119712 264988 119764 264994
rect 119712 264930 119764 264936
rect 106924 264240 106976 264246
rect 106924 264182 106976 264188
rect 116768 264036 116820 264042
rect 116768 263978 116820 263984
rect 112720 263900 112772 263906
rect 112720 263842 112772 263848
rect 3516 263152 3568 263158
rect 3516 263094 3568 263100
rect 3424 262880 3476 262886
rect 3424 262822 3476 262828
rect 2780 215280 2832 215286
rect 2780 215222 2832 215228
rect 2792 214985 2820 215222
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 3436 201929 3464 262822
rect 3528 254153 3556 263094
rect 112536 262812 112588 262818
rect 112536 262754 112588 262760
rect 14464 261316 14516 261322
rect 14464 261258 14516 261264
rect 4804 260364 4856 260370
rect 4804 260306 4856 260312
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 4816 215286 4844 260306
rect 14476 241466 14504 261258
rect 111248 261248 111300 261254
rect 111248 261190 111300 261196
rect 110880 261112 110932 261118
rect 110880 261054 110932 261060
rect 14464 241460 14516 241466
rect 14464 241402 14516 241408
rect 4804 215280 4856 215286
rect 4804 215222 4856 215228
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 107382 200560 107438 200569
rect 107382 200495 107438 200504
rect 108948 200524 109000 200530
rect 107290 200424 107346 200433
rect 107290 200359 107346 200368
rect 106094 199608 106150 199617
rect 106094 199543 106150 199552
rect 102046 199064 102102 199073
rect 102046 198999 102102 199008
rect 100574 197976 100630 197985
rect 100574 197911 100630 197920
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3436 151814 3464 162823
rect 3436 151786 3556 151814
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 149122 3464 149767
rect 3424 149116 3476 149122
rect 3424 149058 3476 149064
rect 3528 145586 3556 151786
rect 9588 149116 9640 149122
rect 9588 149058 9640 149064
rect 9600 148374 9628 149058
rect 100208 148640 100260 148646
rect 100208 148582 100260 148588
rect 9588 148368 9640 148374
rect 9588 148310 9640 148316
rect 3516 145580 3568 145586
rect 3516 145522 3568 145528
rect 3424 142180 3476 142186
rect 3424 142122 3476 142128
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 2780 78056 2832 78062
rect 2780 77998 2832 78004
rect 572 4140 624 4146
rect 572 4082 624 4088
rect 584 480 612 4082
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1688 480 1716 4014
rect 2792 3534 2820 77998
rect 2872 77988 2924 77994
rect 2872 77930 2924 77936
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 77930
rect 3436 45529 3464 142122
rect 17224 141024 17276 141030
rect 17224 140966 17276 140972
rect 8944 140956 8996 140962
rect 8944 140898 8996 140904
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 6920 78124 6972 78130
rect 6920 78066 6972 78072
rect 3516 71664 3568 71670
rect 3514 71632 3516 71641
rect 3568 71632 3570 71641
rect 3514 71567 3570 71576
rect 4160 64184 4212 64190
rect 4160 64126 4212 64132
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 4172 16574 4200 64126
rect 6932 16574 6960 78066
rect 7564 75200 7616 75206
rect 7564 75142 7616 75148
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5276 480 5304 16546
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 7484 3482 7512 16546
rect 7576 4146 7604 75142
rect 8956 71670 8984 140898
rect 14464 72480 14516 72486
rect 14464 72422 14516 72428
rect 8944 71664 8996 71670
rect 8944 71606 8996 71612
rect 8942 68232 8998 68241
rect 8942 68167 8998 68176
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 8956 4078 8984 68167
rect 11058 66872 11114 66881
rect 11058 66807 11114 66816
rect 10324 62824 10376 62830
rect 10324 62766 10376 62772
rect 9680 53100 9732 53106
rect 9680 53042 9732 53048
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 6472 480 6500 3470
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8772 480 8800 3402
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 53042
rect 10336 3466 10364 62766
rect 11072 16574 11100 66807
rect 12440 55888 12492 55894
rect 12440 55830 12492 55836
rect 12452 16574 12480 55830
rect 13820 40724 13872 40730
rect 13820 40666 13872 40672
rect 13832 16574 13860 40666
rect 11072 16546 11192 16574
rect 12452 16546 13584 16574
rect 13832 16546 14320 16574
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11164 480 11192 16546
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12360 480 12388 2926
rect 13556 480 13584 16546
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 14476 2990 14504 72422
rect 17236 6866 17264 140966
rect 31022 139496 31078 139505
rect 31022 139431 31078 139440
rect 31036 111790 31064 139431
rect 31024 111784 31076 111790
rect 31024 111726 31076 111732
rect 95238 81560 95294 81569
rect 95238 81495 95294 81504
rect 71780 80708 71832 80714
rect 71780 80650 71832 80656
rect 57980 78328 58032 78334
rect 57980 78270 58032 78276
rect 46940 78260 46992 78266
rect 46940 78202 46992 78208
rect 20720 78192 20772 78198
rect 20720 78134 20772 78140
rect 18604 69692 18656 69698
rect 18604 69634 18656 69640
rect 17960 60036 18012 60042
rect 17960 59978 18012 59984
rect 17314 36544 17370 36553
rect 17314 36479 17370 36488
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17328 4146 17356 36479
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 15948 480 15976 4082
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17052 480 17080 3402
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 59978
rect 18616 3466 18644 69634
rect 20732 16574 20760 78134
rect 35900 76560 35952 76566
rect 34518 76528 34574 76537
rect 35900 76502 35952 76508
rect 34518 76463 34574 76472
rect 22744 75268 22796 75274
rect 22744 75210 22796 75216
rect 21364 73840 21416 73846
rect 21364 73782 21416 73788
rect 20732 16546 21312 16574
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 19444 480 19472 3538
rect 21284 3482 21312 16546
rect 21376 3602 21404 73782
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21284 3454 21864 3482
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20640 480 20668 2994
rect 21836 480 21864 3454
rect 22756 3058 22784 75210
rect 23480 72548 23532 72554
rect 23480 72490 23532 72496
rect 23492 16574 23520 72490
rect 27620 71188 27672 71194
rect 27620 71130 27672 71136
rect 26240 71120 26292 71126
rect 26240 71062 26292 71068
rect 25502 57216 25558 57225
rect 25502 57151 25558 57160
rect 24858 33824 24914 33833
rect 24858 33759 24914 33768
rect 24872 16574 24900 33759
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23032 480 23060 2994
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 25516 3058 25544 57151
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 71062
rect 27632 3466 27660 71130
rect 27710 51776 27766 51785
rect 27710 51711 27766 51720
rect 27620 3460 27672 3466
rect 27620 3402 27672 3408
rect 27724 480 27752 51711
rect 30378 50280 30434 50289
rect 30378 50215 30434 50224
rect 30392 16574 30420 50215
rect 31760 39364 31812 39370
rect 31760 39306 31812 39312
rect 31772 16574 31800 39306
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 30104 7608 30156 7614
rect 30104 7550 30156 7556
rect 28540 3460 28592 3466
rect 28540 3402 28592 3408
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3402
rect 30116 480 30144 7550
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33612 480 33640 3402
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 76463
rect 35912 6914 35940 76502
rect 45560 71052 45612 71058
rect 45560 70994 45612 71000
rect 41418 69592 41474 69601
rect 41418 69527 41474 69536
rect 40038 67008 40094 67017
rect 40038 66943 40094 66952
rect 35992 65544 36044 65550
rect 35992 65486 36044 65492
rect 36004 16574 36032 65486
rect 39302 48920 39358 48929
rect 39302 48855 39358 48864
rect 38660 37936 38712 37942
rect 38660 37878 38712 37884
rect 38672 16574 38700 37878
rect 36004 16546 36768 16574
rect 38672 16546 39160 16574
rect 35912 6886 36032 6914
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 480 38424 3130
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39316 3194 39344 48855
rect 40052 16574 40080 66943
rect 41432 16574 41460 69527
rect 42800 61396 42852 61402
rect 42800 61338 42852 61344
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 42812 354 42840 61338
rect 44178 47560 44234 47569
rect 44178 47495 44234 47504
rect 44192 3602 44220 47495
rect 44272 31068 44324 31074
rect 44272 31010 44324 31016
rect 44180 3596 44232 3602
rect 44180 3538 44232 3544
rect 44284 480 44312 31010
rect 45572 16574 45600 70994
rect 46204 69760 46256 69766
rect 46204 69702 46256 69708
rect 45572 16546 46152 16574
rect 45928 3936 45980 3942
rect 45928 3878 45980 3884
rect 45100 3596 45152 3602
rect 45100 3538 45152 3544
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45112 354 45140 3538
rect 45940 3466 45968 3878
rect 46124 3482 46152 16546
rect 46216 3942 46244 69702
rect 46952 16574 46980 78202
rect 52460 76628 52512 76634
rect 52460 76570 52512 76576
rect 48320 68332 48372 68338
rect 48320 68274 48372 68280
rect 48332 16574 48360 68274
rect 49700 58676 49752 58682
rect 49700 58618 49752 58624
rect 49712 16574 49740 58618
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 46204 3936 46256 3942
rect 46204 3878 46256 3884
rect 45928 3460 45980 3466
rect 46124 3454 46704 3482
rect 45928 3402 45980 3408
rect 46676 480 46704 3454
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 51356 3596 51408 3602
rect 51356 3538 51408 3544
rect 51368 480 51396 3538
rect 52472 3466 52500 76570
rect 54484 73908 54536 73914
rect 54484 73850 54536 73856
rect 52552 61464 52604 61470
rect 52552 61406 52604 61412
rect 52460 3460 52512 3466
rect 52460 3402 52512 3408
rect 52564 480 52592 61406
rect 53840 35216 53892 35222
rect 53840 35158 53892 35164
rect 53852 16574 53880 35158
rect 53852 16546 54432 16574
rect 54404 3482 54432 16546
rect 54496 3602 54524 73850
rect 57242 65512 57298 65521
rect 57242 65447 57298 65456
rect 56598 46200 56654 46209
rect 56598 46135 56654 46144
rect 56612 16574 56640 46135
rect 56612 16546 56824 16574
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 53380 3460 53432 3466
rect 54404 3454 54984 3482
rect 53380 3402 53432 3408
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3402
rect 54956 480 54984 3454
rect 56048 3460 56100 3466
rect 56048 3402 56100 3408
rect 56060 480 56088 3402
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 57256 3466 57284 65447
rect 57992 16574 58020 78270
rect 60738 77888 60794 77897
rect 60738 77823 60794 77832
rect 57992 16546 58480 16574
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 58452 480 58480 16546
rect 59636 3596 59688 3602
rect 59636 3538 59688 3544
rect 59648 480 59676 3538
rect 60752 3466 60780 77823
rect 64144 76696 64196 76702
rect 64144 76638 64196 76644
rect 62120 64252 62172 64258
rect 62120 64194 62172 64200
rect 60832 44872 60884 44878
rect 60832 44814 60884 44820
rect 60740 3460 60792 3466
rect 60740 3402 60792 3408
rect 60844 480 60872 44814
rect 62132 16574 62160 64194
rect 63500 55956 63552 55962
rect 63500 55898 63552 55904
rect 63512 16574 63540 55898
rect 62132 16546 63264 16574
rect 63512 16546 64092 16574
rect 61660 3460 61712 3466
rect 61660 3402 61712 3408
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61672 354 61700 3402
rect 63236 480 63264 16546
rect 64064 3482 64092 16546
rect 64156 3602 64184 76638
rect 67640 75336 67692 75342
rect 67640 75278 67692 75284
rect 66720 3664 66772 3670
rect 66720 3606 66772 3612
rect 64144 3596 64196 3602
rect 64144 3538 64196 3544
rect 64064 3454 64368 3482
rect 64340 480 64368 3454
rect 65524 3460 65576 3466
rect 65524 3402 65576 3408
rect 65536 480 65564 3402
rect 66732 480 66760 3606
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 75278
rect 70400 72616 70452 72622
rect 70400 72558 70452 72564
rect 69020 60104 69072 60110
rect 69020 60046 69072 60052
rect 69032 16574 69060 60046
rect 70412 16574 70440 72558
rect 71792 16574 71820 80650
rect 72424 76764 72476 76770
rect 72424 76706 72476 76712
rect 69032 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72372 16574
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 69124 480 69152 3538
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72344 3482 72372 16546
rect 72436 3670 72464 76706
rect 81440 75404 81492 75410
rect 81440 75346 81492 75352
rect 78680 68468 78732 68474
rect 78680 68410 78732 68416
rect 75920 68400 75972 68406
rect 75920 68342 75972 68348
rect 75182 62792 75238 62801
rect 75182 62727 75238 62736
rect 74538 43480 74594 43489
rect 74538 43415 74594 43424
rect 74552 16574 74580 43415
rect 74552 16546 75040 16574
rect 73804 4140 73856 4146
rect 73804 4082 73856 4088
rect 72424 3664 72476 3670
rect 72424 3606 72476 3612
rect 72344 3454 72648 3482
rect 72620 480 72648 3454
rect 73816 480 73844 4082
rect 75012 480 75040 16546
rect 75196 4146 75224 62727
rect 75184 4140 75236 4146
rect 75184 4082 75236 4088
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 68342
rect 77298 57352 77354 57361
rect 77298 57287 77354 57296
rect 77312 6914 77340 57287
rect 77392 42084 77444 42090
rect 77392 42026 77444 42032
rect 77404 16574 77432 42026
rect 78692 16574 78720 68410
rect 80060 67040 80112 67046
rect 80060 66982 80112 66988
rect 80072 16574 80100 66982
rect 81452 16574 81480 75346
rect 93860 74044 93912 74050
rect 93860 73986 93912 73992
rect 89720 68604 89772 68610
rect 89720 68546 89772 68552
rect 85580 68536 85632 68542
rect 85580 68478 85632 68484
rect 84198 54496 84254 54505
rect 84198 54431 84254 54440
rect 77404 16546 78168 16574
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 77312 6886 77432 6914
rect 77404 480 77432 6886
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83280 3664 83332 3670
rect 83280 3606 83332 3612
rect 83292 480 83320 3606
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 54431
rect 85592 16574 85620 68478
rect 88340 62892 88392 62898
rect 88340 62834 88392 62840
rect 88352 16574 88380 62834
rect 89732 16574 89760 68546
rect 92480 67176 92532 67182
rect 92480 67118 92532 67124
rect 85592 16546 86448 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 85672 3732 85724 3738
rect 85672 3674 85724 3680
rect 85684 480 85712 3674
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 87512 10328 87564 10334
rect 87512 10270 87564 10276
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 10270
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91560 3800 91612 3806
rect 91560 3742 91612 3748
rect 91572 480 91600 3742
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 67118
rect 93872 6914 93900 73986
rect 93952 67108 94004 67114
rect 93952 67050 94004 67056
rect 93964 16574 93992 67050
rect 95252 16574 95280 81495
rect 96618 75168 96674 75177
rect 96618 75103 96674 75112
rect 96632 16574 96660 75103
rect 100220 74186 100248 148582
rect 100392 148572 100444 148578
rect 100392 148514 100444 148520
rect 100300 148504 100352 148510
rect 100300 148446 100352 148452
rect 100208 74180 100260 74186
rect 100208 74122 100260 74128
rect 100220 73846 100248 74122
rect 100208 73840 100260 73846
rect 100208 73782 100260 73788
rect 100312 72554 100340 148446
rect 100300 72548 100352 72554
rect 100300 72490 100352 72496
rect 100404 71670 100432 148514
rect 100482 148336 100538 148345
rect 100482 148271 100538 148280
rect 99380 71664 99432 71670
rect 99380 71606 99432 71612
rect 100392 71664 100444 71670
rect 100392 71606 100444 71612
rect 99392 71194 99420 71606
rect 99380 71188 99432 71194
rect 99380 71130 99432 71136
rect 99380 66904 99432 66910
rect 99380 66846 99432 66852
rect 98000 65612 98052 65618
rect 98000 65554 98052 65560
rect 98012 16574 98040 65554
rect 99392 16574 99420 66846
rect 99472 60716 99524 60722
rect 99472 60658 99524 60664
rect 99484 60042 99512 60658
rect 99472 60036 99524 60042
rect 99472 59978 99524 59984
rect 99472 56568 99524 56574
rect 99472 56510 99524 56516
rect 99484 55894 99512 56510
rect 99472 55888 99524 55894
rect 99472 55830 99524 55836
rect 100496 53786 100524 148271
rect 100588 60722 100616 197911
rect 100668 195696 100720 195702
rect 100668 195638 100720 195644
rect 100576 60716 100628 60722
rect 100576 60658 100628 60664
rect 100680 56574 100708 195638
rect 101680 195492 101732 195498
rect 101680 195434 101732 195440
rect 101588 190052 101640 190058
rect 101588 189994 101640 190000
rect 101600 77217 101628 189994
rect 100758 77208 100814 77217
rect 100758 77143 100814 77152
rect 101586 77208 101642 77217
rect 101586 77143 101642 77152
rect 100772 76537 100800 77143
rect 100758 76528 100814 76537
rect 100758 76463 100814 76472
rect 101692 57905 101720 195434
rect 101864 192976 101916 192982
rect 101864 192918 101916 192924
rect 101772 189848 101824 189854
rect 101772 189790 101824 189796
rect 100758 57896 100814 57905
rect 100758 57831 100814 57840
rect 101678 57896 101734 57905
rect 101678 57831 101734 57840
rect 100772 57225 100800 57831
rect 100758 57216 100814 57225
rect 100758 57151 100814 57160
rect 100668 56568 100720 56574
rect 100668 56510 100720 56516
rect 100484 53780 100536 53786
rect 100484 53722 100536 53728
rect 100496 53106 100524 53722
rect 100484 53100 100536 53106
rect 100484 53042 100536 53048
rect 100758 52456 100814 52465
rect 100758 52391 100814 52400
rect 100772 51785 100800 52391
rect 100758 51776 100814 51785
rect 100758 51711 100814 51720
rect 100760 51060 100812 51066
rect 100760 51002 100812 51008
rect 93964 16546 94728 16574
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 93872 6886 93992 6914
rect 93964 480 93992 6886
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 51002
rect 100850 50960 100906 50969
rect 100850 50895 100906 50904
rect 100864 50289 100892 50895
rect 100850 50280 100906 50289
rect 100850 50215 100906 50224
rect 101784 49609 101812 189790
rect 101876 50969 101904 192918
rect 101956 189916 102008 189922
rect 101956 189858 102008 189864
rect 101862 50960 101918 50969
rect 101862 50895 101918 50904
rect 100850 49600 100906 49609
rect 100850 49535 100906 49544
rect 101770 49600 101826 49609
rect 101770 49535 101826 49544
rect 100864 48929 100892 49535
rect 100850 48920 100906 48929
rect 100850 48855 100906 48864
rect 101968 48249 101996 189858
rect 102060 52465 102088 198999
rect 104440 198212 104492 198218
rect 104440 198154 104492 198160
rect 103060 198144 103112 198150
rect 103060 198086 103112 198092
rect 102784 198008 102836 198014
rect 102784 197950 102836 197956
rect 102796 78606 102824 197950
rect 102968 194132 103020 194138
rect 102968 194074 103020 194080
rect 102876 190120 102928 190126
rect 102876 190062 102928 190068
rect 102140 78600 102192 78606
rect 102140 78542 102192 78548
rect 102784 78600 102836 78606
rect 102784 78542 102836 78548
rect 102152 78198 102180 78542
rect 102140 78192 102192 78198
rect 102140 78134 102192 78140
rect 102140 71120 102192 71126
rect 102140 71062 102192 71068
rect 102152 70854 102180 71062
rect 102140 70848 102192 70854
rect 102140 70790 102192 70796
rect 102888 69601 102916 190062
rect 102980 69766 103008 194074
rect 103072 70854 103100 198086
rect 103152 198076 103204 198082
rect 103152 198018 103204 198024
rect 103060 70848 103112 70854
rect 103060 70790 103112 70796
rect 102968 69760 103020 69766
rect 102968 69702 103020 69708
rect 103164 69630 103192 198018
rect 104254 197024 104310 197033
rect 104254 196959 104310 196968
rect 103244 194404 103296 194410
rect 103244 194346 103296 194352
rect 103152 69624 103204 69630
rect 102874 69592 102930 69601
rect 103152 69566 103204 69572
rect 102874 69527 102930 69536
rect 102140 66972 102192 66978
rect 102140 66914 102192 66920
rect 102046 52456 102102 52465
rect 102046 52391 102102 52400
rect 100850 48240 100906 48249
rect 100850 48175 100906 48184
rect 101954 48240 102010 48249
rect 101954 48175 102010 48184
rect 100864 47569 100892 48175
rect 100850 47560 100906 47569
rect 100850 47495 100906 47504
rect 102152 3398 102180 66914
rect 103256 66230 103284 194346
rect 104164 194200 104216 194206
rect 104164 194142 104216 194148
rect 103428 193996 103480 194002
rect 103428 193938 103480 193944
rect 103336 193928 103388 193934
rect 103336 193870 103388 193876
rect 102232 66224 102284 66230
rect 102232 66166 102284 66172
rect 103244 66224 103296 66230
rect 103244 66166 103296 66172
rect 102244 65550 102272 66166
rect 102232 65544 102284 65550
rect 102232 65486 102284 65492
rect 103348 64870 103376 193870
rect 102232 64864 102284 64870
rect 102232 64806 102284 64812
rect 103336 64864 103388 64870
rect 103336 64806 103388 64812
rect 102244 64258 102272 64806
rect 102232 64252 102284 64258
rect 102232 64194 102284 64200
rect 103440 62082 103468 193938
rect 104072 193724 104124 193730
rect 104072 193666 104124 193672
rect 104084 78470 104112 193666
rect 104072 78464 104124 78470
rect 104072 78406 104124 78412
rect 104084 78062 104112 78406
rect 104072 78056 104124 78062
rect 104072 77998 104124 78004
rect 104176 74118 104204 194142
rect 104164 74112 104216 74118
rect 104164 74054 104216 74060
rect 104268 73982 104296 196959
rect 104348 191140 104400 191146
rect 104348 191082 104400 191088
rect 104256 73976 104308 73982
rect 104256 73918 104308 73924
rect 104256 73364 104308 73370
rect 104256 73306 104308 73312
rect 103520 69556 103572 69562
rect 103520 69498 103572 69504
rect 102232 62076 102284 62082
rect 102232 62018 102284 62024
rect 103428 62076 103480 62082
rect 103428 62018 103480 62024
rect 102244 61470 102272 62018
rect 102232 61464 102284 61470
rect 102232 61406 102284 61412
rect 102232 53100 102284 53106
rect 102232 53042 102284 53048
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 53042
rect 103532 16574 103560 69498
rect 104268 67561 104296 73306
rect 104360 67590 104388 191082
rect 104452 72758 104480 198154
rect 106004 196784 106056 196790
rect 106004 196726 106056 196732
rect 105728 195424 105780 195430
rect 105728 195366 105780 195372
rect 104532 194336 104584 194342
rect 104532 194278 104584 194284
rect 104440 72752 104492 72758
rect 104440 72694 104492 72700
rect 104452 72486 104480 72694
rect 104440 72480 104492 72486
rect 104440 72422 104492 72428
rect 104544 70530 104572 194278
rect 104624 194268 104676 194274
rect 104624 194210 104676 194216
rect 104636 73370 104664 194210
rect 104714 193896 104770 193905
rect 104714 193831 104770 193840
rect 104624 73364 104676 73370
rect 104624 73306 104676 73312
rect 104544 70502 104664 70530
rect 104636 68814 104664 70502
rect 104624 68808 104676 68814
rect 104624 68750 104676 68756
rect 104636 68338 104664 68750
rect 104624 68332 104676 68338
rect 104624 68274 104676 68280
rect 104348 67584 104400 67590
rect 104254 67552 104310 67561
rect 104348 67526 104400 67532
rect 104254 67487 104310 67496
rect 104360 67046 104388 67526
rect 104348 67040 104400 67046
rect 104348 66982 104400 66988
rect 104728 63510 104756 193831
rect 104808 191208 104860 191214
rect 104808 191150 104860 191156
rect 104716 63504 104768 63510
rect 104716 63446 104768 63452
rect 104728 62830 104756 63446
rect 104716 62824 104768 62830
rect 104716 62766 104768 62772
rect 104820 60654 104848 191150
rect 105636 148436 105688 148442
rect 105636 148378 105688 148384
rect 104900 79348 104952 79354
rect 104900 79290 104952 79296
rect 104912 75886 104940 79290
rect 105544 77240 105596 77246
rect 105544 77182 105596 77188
rect 105556 76362 105584 77182
rect 105544 76356 105596 76362
rect 105544 76298 105596 76304
rect 104900 75880 104952 75886
rect 104900 75822 104952 75828
rect 104912 74050 104940 75822
rect 104900 74044 104952 74050
rect 104900 73986 104952 73992
rect 105450 66192 105506 66201
rect 105450 66127 105506 66136
rect 105464 65521 105492 66127
rect 105450 65512 105506 65521
rect 105450 65447 105506 65456
rect 104808 60648 104860 60654
rect 104808 60590 104860 60596
rect 104820 60110 104848 60590
rect 104808 60104 104860 60110
rect 104808 60046 104860 60052
rect 105556 51066 105584 76298
rect 105648 73001 105676 148378
rect 105740 80209 105768 195366
rect 105912 194472 105964 194478
rect 105912 194414 105964 194420
rect 105820 193860 105872 193866
rect 105820 193802 105872 193808
rect 105726 80200 105782 80209
rect 105726 80135 105782 80144
rect 105634 72992 105690 73001
rect 105634 72927 105690 72936
rect 105648 67182 105676 72927
rect 105740 68610 105768 80135
rect 105832 77246 105860 193802
rect 105924 79234 105952 194414
rect 106016 79354 106044 196726
rect 106004 79348 106056 79354
rect 106004 79290 106056 79296
rect 105924 79206 106044 79234
rect 105820 77240 105872 77246
rect 105820 77182 105872 77188
rect 106016 76974 106044 79206
rect 106004 76968 106056 76974
rect 106004 76910 106056 76916
rect 106016 76702 106044 76910
rect 106004 76696 106056 76702
rect 106004 76638 106056 76644
rect 106108 72962 106136 199543
rect 107108 198416 107160 198422
rect 107108 198358 107160 198364
rect 106188 194540 106240 194546
rect 106188 194482 106240 194488
rect 106096 72956 106148 72962
rect 106096 72898 106148 72904
rect 105728 68604 105780 68610
rect 105728 68546 105780 68552
rect 106108 68542 106136 72898
rect 106096 68536 106148 68542
rect 106096 68478 106148 68484
rect 105636 67176 105688 67182
rect 105636 67118 105688 67124
rect 106200 66201 106228 194482
rect 107016 194064 107068 194070
rect 107016 194006 107068 194012
rect 106924 193792 106976 193798
rect 106924 193734 106976 193740
rect 106832 189780 106884 189786
rect 106832 189722 106884 189728
rect 106740 80436 106792 80442
rect 106740 80378 106792 80384
rect 106752 75721 106780 80378
rect 106844 79490 106872 189722
rect 106832 79484 106884 79490
rect 106832 79426 106884 79432
rect 106936 76838 106964 193734
rect 107028 80442 107056 194006
rect 107016 80436 107068 80442
rect 107016 80378 107068 80384
rect 107016 80300 107068 80306
rect 107016 80242 107068 80248
rect 106924 76832 106976 76838
rect 106924 76774 106976 76780
rect 107028 75818 107056 80242
rect 107120 78130 107148 198358
rect 107200 197056 107252 197062
rect 107200 196998 107252 197004
rect 107212 80306 107240 196998
rect 107304 89146 107332 200359
rect 107292 89140 107344 89146
rect 107292 89082 107344 89088
rect 107396 89026 107424 200495
rect 108948 200466 109000 200472
rect 107566 198792 107622 198801
rect 107566 198727 107622 198736
rect 107474 196888 107530 196897
rect 107474 196823 107530 196832
rect 107304 88998 107424 89026
rect 107200 80300 107252 80306
rect 107200 80242 107252 80248
rect 107304 80186 107332 88998
rect 107384 88936 107436 88942
rect 107384 88878 107436 88884
rect 107212 80158 107332 80186
rect 107212 78266 107240 80158
rect 107396 80050 107424 88878
rect 107304 80022 107424 80050
rect 107304 78334 107332 80022
rect 107292 78328 107344 78334
rect 107292 78270 107344 78276
rect 107200 78260 107252 78266
rect 107200 78202 107252 78208
rect 107108 78124 107160 78130
rect 107108 78066 107160 78072
rect 107212 77518 107240 78202
rect 107304 77722 107332 78270
rect 107384 78124 107436 78130
rect 107384 78066 107436 78072
rect 107396 77858 107424 78066
rect 107384 77852 107436 77858
rect 107384 77794 107436 77800
rect 107292 77716 107344 77722
rect 107292 77658 107344 77664
rect 107200 77512 107252 77518
rect 107200 77454 107252 77460
rect 107016 75812 107068 75818
rect 107016 75754 107068 75760
rect 106738 75712 106794 75721
rect 106738 75647 106794 75656
rect 107028 68406 107056 75754
rect 107488 72894 107516 196823
rect 107580 73914 107608 198727
rect 108580 198552 108632 198558
rect 108580 198494 108632 198500
rect 108396 197192 108448 197198
rect 108396 197134 108448 197140
rect 108302 192536 108358 192545
rect 108302 192471 108358 192480
rect 108120 189984 108172 189990
rect 108120 189926 108172 189932
rect 108132 142866 108160 189926
rect 108212 148776 108264 148782
rect 108212 148718 108264 148724
rect 108120 142860 108172 142866
rect 108120 142802 108172 142808
rect 107568 73908 107620 73914
rect 107568 73850 107620 73856
rect 107580 73710 107608 73850
rect 107568 73704 107620 73710
rect 107568 73646 107620 73652
rect 107476 72888 107528 72894
rect 107476 72830 107528 72836
rect 107488 68474 107516 72830
rect 107660 70440 107712 70446
rect 107660 70382 107712 70388
rect 107476 68468 107528 68474
rect 107476 68410 107528 68416
rect 107016 68400 107068 68406
rect 107016 68342 107068 68348
rect 106280 67040 106332 67046
rect 106280 66982 106332 66988
rect 106186 66192 106242 66201
rect 106186 66127 106242 66136
rect 105544 51060 105596 51066
rect 105544 51002 105596 51008
rect 106292 16574 106320 66982
rect 107672 16574 107700 70382
rect 108224 55214 108252 148718
rect 108316 80918 108344 192471
rect 108304 80912 108356 80918
rect 108304 80854 108356 80860
rect 108408 80714 108436 197134
rect 108488 195764 108540 195770
rect 108488 195706 108540 195712
rect 108396 80708 108448 80714
rect 108396 80650 108448 80656
rect 108500 77042 108528 195706
rect 108592 77994 108620 198494
rect 108672 198348 108724 198354
rect 108672 198290 108724 198296
rect 108580 77988 108632 77994
rect 108580 77930 108632 77936
rect 108488 77036 108540 77042
rect 108488 76978 108540 76984
rect 108500 69562 108528 76978
rect 108684 75614 108712 198290
rect 108764 195832 108816 195838
rect 108764 195774 108816 195780
rect 108672 75608 108724 75614
rect 108672 75550 108724 75556
rect 108776 71466 108804 195774
rect 108856 192636 108908 192642
rect 108856 192578 108908 192584
rect 108764 71460 108816 71466
rect 108764 71402 108816 71408
rect 108776 70446 108804 71402
rect 108764 70440 108816 70446
rect 108764 70382 108816 70388
rect 108488 69556 108540 69562
rect 108488 69498 108540 69504
rect 108868 68882 108896 192578
rect 108960 71194 108988 200466
rect 110236 196852 110288 196858
rect 110236 196794 110288 196800
rect 110052 196716 110104 196722
rect 110052 196658 110104 196664
rect 109960 196648 110012 196654
rect 109960 196590 110012 196596
rect 109776 192772 109828 192778
rect 109776 192714 109828 192720
rect 109788 79354 109816 192714
rect 109868 192568 109920 192574
rect 109868 192510 109920 192516
rect 109880 79762 109908 192510
rect 109868 79756 109920 79762
rect 109868 79698 109920 79704
rect 109776 79348 109828 79354
rect 109776 79290 109828 79296
rect 109972 74526 110000 196590
rect 109960 74520 110012 74526
rect 109960 74462 110012 74468
rect 110064 74458 110092 196658
rect 110144 190188 110196 190194
rect 110144 190130 110196 190136
rect 110052 74452 110104 74458
rect 110052 74394 110104 74400
rect 108948 71188 109000 71194
rect 108948 71130 109000 71136
rect 109040 69012 109092 69018
rect 109040 68954 109092 68960
rect 108856 68876 108908 68882
rect 108856 68818 108908 68824
rect 108224 55186 108436 55214
rect 108408 44169 108436 55186
rect 108394 44160 108450 44169
rect 108394 44095 108450 44104
rect 108408 43489 108436 44095
rect 108394 43480 108450 43489
rect 108394 43415 108450 43424
rect 103532 16546 104112 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105728 8968 105780 8974
rect 105728 8910 105780 8916
rect 105740 480 105768 8910
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109052 354 109080 68954
rect 110156 67454 110184 190130
rect 110248 73166 110276 196794
rect 110328 191276 110380 191282
rect 110328 191218 110380 191224
rect 110236 73160 110288 73166
rect 110236 73102 110288 73108
rect 110144 67448 110196 67454
rect 110144 67390 110196 67396
rect 110340 57361 110368 191218
rect 110892 147150 110920 261054
rect 111064 261044 111116 261050
rect 111064 260986 111116 260992
rect 110970 189680 111026 189689
rect 110970 189615 111026 189624
rect 110880 147144 110932 147150
rect 110880 147086 110932 147092
rect 110880 147008 110932 147014
rect 110880 146950 110932 146956
rect 110788 144696 110840 144702
rect 110788 144638 110840 144644
rect 110800 75886 110828 144638
rect 110788 75880 110840 75886
rect 110788 75822 110840 75828
rect 110418 63472 110474 63481
rect 110418 63407 110474 63416
rect 110432 62801 110460 63407
rect 110418 62792 110474 62801
rect 110418 62727 110474 62736
rect 110420 59356 110472 59362
rect 110420 59298 110472 59304
rect 110326 57352 110382 57361
rect 110326 57287 110382 57296
rect 110432 16574 110460 59298
rect 110892 46889 110920 146950
rect 110984 75585 111012 189615
rect 111076 144294 111104 260986
rect 111156 196988 111208 196994
rect 111156 196930 111208 196936
rect 111064 144288 111116 144294
rect 111064 144230 111116 144236
rect 111168 79422 111196 196930
rect 111260 142934 111288 261190
rect 111616 200592 111668 200598
rect 111616 200534 111668 200540
rect 111524 195628 111576 195634
rect 111524 195570 111576 195576
rect 111432 192840 111484 192846
rect 111432 192782 111484 192788
rect 111338 192672 111394 192681
rect 111338 192607 111394 192616
rect 111248 142928 111300 142934
rect 111248 142870 111300 142876
rect 111156 79416 111208 79422
rect 111156 79358 111208 79364
rect 111064 75880 111116 75886
rect 111064 75822 111116 75828
rect 111076 75682 111104 75822
rect 111064 75676 111116 75682
rect 111064 75618 111116 75624
rect 110970 75576 111026 75585
rect 110970 75511 111026 75520
rect 110984 69018 111012 75511
rect 110972 69012 111024 69018
rect 110972 68954 111024 68960
rect 111076 65618 111104 75618
rect 111352 73234 111380 192607
rect 111444 74254 111472 192782
rect 111536 74322 111564 195570
rect 111524 74316 111576 74322
rect 111524 74258 111576 74264
rect 111432 74248 111484 74254
rect 111432 74190 111484 74196
rect 111340 73228 111392 73234
rect 111340 73170 111392 73176
rect 111628 72826 111656 200534
rect 112350 192808 112406 192817
rect 112350 192743 112406 192752
rect 111708 191344 111760 191350
rect 111708 191286 111760 191292
rect 111616 72820 111668 72826
rect 111616 72762 111668 72768
rect 111064 65612 111116 65618
rect 111064 65554 111116 65560
rect 111720 63481 111748 191286
rect 112260 148164 112312 148170
rect 112260 148106 112312 148112
rect 111706 63472 111762 63481
rect 111706 63407 111762 63416
rect 112272 59294 112300 148106
rect 112364 79626 112392 192743
rect 112444 192500 112496 192506
rect 112444 192442 112496 192448
rect 112352 79620 112404 79626
rect 112352 79562 112404 79568
rect 112456 76430 112484 192442
rect 112548 146062 112576 262754
rect 112628 260024 112680 260030
rect 112628 259966 112680 259972
rect 112536 146056 112588 146062
rect 112536 145998 112588 146004
rect 112536 145920 112588 145926
rect 112536 145862 112588 145868
rect 112444 76424 112496 76430
rect 112444 76366 112496 76372
rect 112548 74089 112576 145862
rect 112640 142730 112668 259966
rect 112732 146130 112760 263842
rect 114008 263696 114060 263702
rect 114008 263638 114060 263644
rect 113732 262744 113784 262750
rect 113732 262686 113784 262692
rect 112996 195968 113048 195974
rect 112996 195910 113048 195916
rect 112812 195900 112864 195906
rect 112812 195842 112864 195848
rect 112720 146124 112772 146130
rect 112720 146066 112772 146072
rect 112720 144764 112772 144770
rect 112720 144706 112772 144712
rect 112628 142724 112680 142730
rect 112628 142666 112680 142672
rect 112534 74080 112590 74089
rect 112534 74015 112590 74024
rect 112548 67114 112576 74015
rect 112732 69902 112760 144706
rect 112824 73914 112852 195842
rect 112904 195560 112956 195566
rect 112904 195502 112956 195508
rect 112916 74390 112944 195502
rect 112904 74384 112956 74390
rect 112904 74326 112956 74332
rect 112812 73908 112864 73914
rect 112812 73850 112864 73856
rect 113008 73846 113036 195910
rect 113088 191412 113140 191418
rect 113088 191354 113140 191360
rect 112996 73840 113048 73846
rect 112996 73782 113048 73788
rect 112720 69896 112772 69902
rect 112720 69838 112772 69844
rect 112536 67108 112588 67114
rect 112536 67050 112588 67056
rect 111800 59288 111852 59294
rect 111800 59230 111852 59236
rect 112260 59288 112312 59294
rect 112260 59230 112312 59236
rect 111812 58682 111840 59230
rect 111800 58676 111852 58682
rect 111800 58618 111852 58624
rect 113100 55185 113128 191354
rect 113548 148980 113600 148986
rect 113548 148922 113600 148928
rect 113456 146260 113508 146266
rect 113456 146202 113508 146208
rect 113468 71126 113496 146202
rect 113456 71120 113508 71126
rect 113456 71062 113508 71068
rect 113180 68332 113232 68338
rect 113180 68274 113232 68280
rect 111798 55176 111854 55185
rect 111798 55111 111854 55120
rect 113086 55176 113142 55185
rect 113086 55111 113142 55120
rect 111812 54505 111840 55111
rect 111798 54496 111854 54505
rect 111798 54431 111854 54440
rect 110510 46880 110566 46889
rect 110510 46815 110566 46824
rect 110878 46880 110934 46889
rect 110878 46815 110934 46824
rect 110524 46209 110552 46815
rect 110510 46200 110566 46209
rect 110510 46135 110566 46144
rect 113192 16574 113220 68274
rect 113468 64874 113496 71062
rect 113560 69970 113588 148922
rect 113744 145994 113772 262686
rect 113916 262540 113968 262546
rect 113916 262482 113968 262488
rect 113824 197328 113876 197334
rect 113824 197270 113876 197276
rect 113732 145988 113784 145994
rect 113732 145930 113784 145936
rect 113640 140616 113692 140622
rect 113640 140558 113692 140564
rect 113652 78062 113680 140558
rect 113730 138952 113786 138961
rect 113730 138887 113786 138896
rect 113640 78056 113692 78062
rect 113640 77998 113692 78004
rect 113744 76673 113772 138887
rect 113836 79558 113864 197270
rect 113928 144498 113956 262482
rect 114020 144634 114048 263638
rect 116676 262948 116728 262954
rect 116676 262890 116728 262896
rect 116584 262676 116636 262682
rect 116584 262618 116636 262624
rect 116492 262608 116544 262614
rect 116492 262550 116544 262556
rect 114100 260908 114152 260914
rect 114100 260850 114152 260856
rect 114008 144628 114060 144634
rect 114008 144570 114060 144576
rect 113916 144492 113968 144498
rect 113916 144434 113968 144440
rect 114008 143472 114060 143478
rect 114008 143414 114060 143420
rect 113824 79552 113876 79558
rect 113824 79494 113876 79500
rect 113730 76664 113786 76673
rect 113730 76599 113786 76608
rect 113548 69964 113600 69970
rect 113548 69906 113600 69912
rect 114020 67522 114048 143414
rect 114112 141778 114140 260850
rect 115296 259684 115348 259690
rect 115296 259626 115348 259632
rect 114192 197260 114244 197266
rect 114192 197202 114244 197208
rect 114100 141772 114152 141778
rect 114100 141714 114152 141720
rect 114204 73778 114232 197202
rect 114468 197124 114520 197130
rect 114468 197066 114520 197072
rect 114282 195392 114338 195401
rect 114282 195327 114338 195336
rect 114192 73772 114244 73778
rect 114192 73714 114244 73720
rect 114296 70922 114324 195327
rect 114376 193112 114428 193118
rect 114376 193054 114428 193060
rect 114284 70916 114336 70922
rect 114284 70858 114336 70864
rect 114388 68921 114416 193054
rect 114480 71369 114508 197066
rect 114836 192432 114888 192438
rect 114836 192374 114888 192380
rect 114560 73228 114612 73234
rect 114560 73170 114612 73176
rect 114466 71360 114522 71369
rect 114466 71295 114522 71304
rect 114374 68912 114430 68921
rect 114374 68847 114430 68856
rect 114008 67516 114060 67522
rect 114008 67458 114060 67464
rect 113468 64846 113864 64874
rect 113836 53106 113864 64846
rect 113824 53100 113876 53106
rect 113824 53042 113876 53048
rect 114572 16574 114600 73170
rect 114848 68785 114876 192374
rect 115020 149048 115072 149054
rect 115020 148990 115072 148996
rect 114928 148232 114980 148238
rect 114928 148174 114980 148180
rect 114940 73953 114968 148174
rect 114926 73944 114982 73953
rect 114926 73879 114982 73888
rect 114834 68776 114890 68785
rect 114834 68711 114890 68720
rect 114940 64874 114968 73879
rect 115032 69834 115060 148990
rect 115204 147212 115256 147218
rect 115204 147154 115256 147160
rect 115110 139088 115166 139097
rect 115110 139023 115166 139032
rect 115124 70009 115152 139023
rect 115216 75546 115244 147154
rect 115308 146198 115336 259626
rect 115480 259548 115532 259554
rect 115480 259490 115532 259496
rect 115388 193044 115440 193050
rect 115388 192986 115440 192992
rect 115296 146192 115348 146198
rect 115296 146134 115348 146140
rect 115400 75750 115428 192986
rect 115492 141846 115520 259490
rect 115664 199504 115716 199510
rect 115664 199446 115716 199452
rect 115572 191480 115624 191486
rect 115572 191422 115624 191428
rect 115480 141840 115532 141846
rect 115480 141782 115532 141788
rect 115388 75744 115440 75750
rect 115388 75686 115440 75692
rect 115204 75540 115256 75546
rect 115204 75482 115256 75488
rect 115110 70000 115166 70009
rect 115110 69935 115166 69944
rect 115020 69828 115072 69834
rect 115020 69770 115072 69776
rect 115584 69766 115612 191422
rect 115676 77081 115704 199446
rect 115756 199436 115808 199442
rect 115756 199378 115808 199384
rect 115662 77072 115718 77081
rect 115662 77007 115718 77016
rect 115768 75041 115796 199378
rect 116216 145648 116268 145654
rect 116216 145590 116268 145596
rect 116228 79694 116256 145590
rect 116306 144664 116362 144673
rect 116306 144599 116362 144608
rect 116216 79688 116268 79694
rect 116216 79630 116268 79636
rect 115754 75032 115810 75041
rect 115754 74967 115810 74976
rect 115848 73228 115900 73234
rect 115848 73170 115900 73176
rect 115860 72690 115888 73170
rect 115848 72684 115900 72690
rect 115848 72626 115900 72632
rect 115940 71800 115992 71806
rect 116320 71777 116348 144599
rect 116504 144566 116532 262550
rect 116492 144560 116544 144566
rect 116492 144502 116544 144508
rect 116596 143342 116624 262618
rect 116688 143546 116716 262890
rect 116676 143540 116728 143546
rect 116676 143482 116728 143488
rect 116584 143336 116636 143342
rect 116584 143278 116636 143284
rect 116780 143274 116808 263978
rect 119528 263968 119580 263974
rect 119528 263910 119580 263916
rect 118424 262472 118476 262478
rect 118424 262414 118476 262420
rect 118240 262404 118292 262410
rect 118240 262346 118292 262352
rect 116860 262268 116912 262274
rect 116860 262210 116912 262216
rect 116768 143268 116820 143274
rect 116768 143210 116820 143216
rect 116492 142860 116544 142866
rect 116492 142802 116544 142808
rect 116400 140344 116452 140350
rect 116400 140286 116452 140292
rect 116412 80753 116440 140286
rect 116398 80744 116454 80753
rect 116398 80679 116454 80688
rect 116504 72486 116532 142802
rect 116872 141302 116900 262210
rect 117964 261180 118016 261186
rect 117964 261122 118016 261128
rect 117872 259616 117924 259622
rect 117872 259558 117924 259564
rect 117044 199572 117096 199578
rect 117044 199514 117096 199520
rect 116952 192908 117004 192914
rect 116952 192850 117004 192856
rect 116860 141296 116912 141302
rect 116860 141238 116912 141244
rect 116584 140276 116636 140282
rect 116584 140218 116636 140224
rect 116596 80714 116624 140218
rect 116768 140140 116820 140146
rect 116768 140082 116820 140088
rect 116584 80708 116636 80714
rect 116584 80650 116636 80656
rect 116492 72480 116544 72486
rect 116492 72422 116544 72428
rect 116504 71806 116532 72422
rect 116492 71800 116544 71806
rect 115940 71742 115992 71748
rect 116306 71768 116362 71777
rect 115572 69760 115624 69766
rect 115572 69702 115624 69708
rect 114940 64846 115244 64874
rect 115216 59362 115244 64846
rect 115204 59356 115256 59362
rect 115204 59298 115256 59304
rect 115952 16574 115980 71742
rect 116492 71742 116544 71748
rect 116306 71703 116362 71712
rect 116780 71505 116808 140082
rect 116964 71534 116992 192850
rect 117056 76945 117084 199514
rect 117136 196920 117188 196926
rect 117136 196862 117188 196868
rect 117042 76936 117098 76945
rect 117042 76871 117098 76880
rect 117148 72729 117176 196862
rect 117228 192704 117280 192710
rect 117228 192646 117280 192652
rect 117134 72720 117190 72729
rect 117134 72655 117190 72664
rect 116952 71528 117004 71534
rect 116766 71496 116822 71505
rect 116952 71470 117004 71476
rect 116766 71431 116822 71440
rect 117240 68950 117268 192646
rect 117884 189038 117912 259558
rect 117872 189032 117924 189038
rect 117872 188974 117924 188980
rect 117976 147286 118004 261122
rect 118148 259956 118200 259962
rect 118148 259898 118200 259904
rect 118056 259820 118108 259826
rect 118056 259762 118108 259768
rect 117964 147280 118016 147286
rect 117964 147222 118016 147228
rect 118068 147098 118096 259762
rect 117688 147076 117740 147082
rect 117688 147018 117740 147024
rect 117884 147070 118096 147098
rect 117596 146940 117648 146946
rect 117596 146882 117648 146888
rect 117504 145784 117556 145790
rect 117504 145726 117556 145732
rect 117412 76696 117464 76702
rect 117412 76638 117464 76644
rect 117424 75546 117452 76638
rect 117412 75540 117464 75546
rect 117412 75482 117464 75488
rect 117228 68944 117280 68950
rect 117228 68886 117280 68892
rect 117320 68400 117372 68406
rect 117320 68342 117372 68348
rect 110432 16546 110552 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 110524 480 110552 16546
rect 112812 3868 112864 3874
rect 112812 3810 112864 3816
rect 111614 3360 111670 3369
rect 111614 3295 111670 3304
rect 111628 480 111656 3295
rect 112824 480 112852 3810
rect 114020 480 114048 16546
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 68342
rect 117424 3874 117452 75482
rect 117516 71602 117544 145726
rect 117608 78946 117636 146882
rect 117596 78940 117648 78946
rect 117596 78882 117648 78888
rect 117504 71596 117556 71602
rect 117504 71538 117556 71544
rect 117700 70990 117728 147018
rect 117884 144362 117912 147070
rect 117962 146976 118018 146985
rect 117962 146911 118018 146920
rect 117872 144356 117924 144362
rect 117872 144298 117924 144304
rect 117976 141982 118004 146911
rect 118160 143206 118188 259898
rect 118252 144226 118280 262346
rect 118332 261384 118384 261390
rect 118332 261326 118384 261332
rect 118344 146826 118372 261326
rect 118436 146985 118464 262414
rect 119344 259888 119396 259894
rect 119344 259830 119396 259836
rect 118516 199640 118568 199646
rect 118516 199582 118568 199588
rect 118422 146976 118478 146985
rect 118422 146911 118478 146920
rect 118344 146798 118464 146826
rect 118330 144800 118386 144809
rect 118330 144735 118386 144744
rect 118240 144220 118292 144226
rect 118240 144162 118292 144168
rect 118344 143614 118372 144735
rect 118332 143608 118384 143614
rect 118332 143550 118384 143556
rect 118436 143410 118464 146798
rect 118424 143404 118476 143410
rect 118424 143346 118476 143352
rect 118148 143200 118200 143206
rect 118148 143142 118200 143148
rect 118332 142792 118384 142798
rect 118332 142734 118384 142740
rect 117964 141976 118016 141982
rect 117964 141918 118016 141924
rect 118148 141636 118200 141642
rect 118148 141578 118200 141584
rect 117964 141092 118016 141098
rect 117964 141034 118016 141040
rect 117872 140208 117924 140214
rect 117872 140150 117924 140156
rect 117884 78878 117912 140150
rect 117976 137970 118004 141034
rect 118056 139732 118108 139738
rect 118056 139674 118108 139680
rect 117964 137964 118016 137970
rect 117964 137906 118016 137912
rect 118068 136082 118096 139674
rect 117976 136054 118096 136082
rect 117976 79529 118004 136054
rect 118160 122834 118188 141578
rect 118068 122806 118188 122834
rect 117962 79520 118018 79529
rect 117962 79455 118018 79464
rect 118068 79014 118096 122806
rect 118056 79008 118108 79014
rect 118056 78950 118108 78956
rect 117872 78872 117924 78878
rect 117872 78814 117924 78820
rect 117688 70984 117740 70990
rect 117688 70926 117740 70932
rect 118344 69018 118372 142734
rect 118528 76906 118556 199582
rect 118606 196752 118662 196761
rect 118606 196687 118662 196696
rect 118516 76900 118568 76906
rect 118516 76842 118568 76848
rect 118620 72865 118648 196687
rect 119068 145852 119120 145858
rect 119068 145794 119120 145800
rect 118976 145716 119028 145722
rect 118976 145658 119028 145664
rect 118988 77110 119016 145658
rect 118976 77104 119028 77110
rect 118976 77046 119028 77052
rect 118606 72856 118662 72865
rect 118606 72791 118662 72800
rect 119080 71330 119108 145794
rect 119356 142769 119384 259830
rect 119436 259752 119488 259758
rect 119436 259694 119488 259700
rect 119342 142760 119398 142769
rect 119342 142695 119398 142704
rect 119448 141438 119476 259694
rect 119540 143070 119568 263910
rect 119620 263764 119672 263770
rect 119620 263706 119672 263712
rect 119528 143064 119580 143070
rect 119528 143006 119580 143012
rect 119632 143002 119660 263706
rect 119724 144430 119752 264930
rect 119896 264104 119948 264110
rect 119896 264046 119948 264052
rect 119804 260772 119856 260778
rect 119804 260714 119856 260720
rect 119712 144424 119764 144430
rect 119712 144366 119764 144372
rect 119620 142996 119672 143002
rect 119620 142938 119672 142944
rect 119436 141432 119488 141438
rect 119436 141374 119488 141380
rect 119816 141370 119844 260714
rect 119908 141710 119936 264046
rect 133156 263906 133184 271866
rect 134432 264036 134484 264042
rect 134432 263978 134484 263984
rect 133144 263900 133196 263906
rect 133144 263842 133196 263848
rect 120908 263832 120960 263838
rect 120908 263774 120960 263780
rect 120816 260840 120868 260846
rect 120816 260782 120868 260788
rect 120724 259480 120776 259486
rect 120724 259422 120776 259428
rect 119986 200696 120042 200705
rect 119986 200631 120042 200640
rect 119896 141704 119948 141710
rect 119896 141646 119948 141652
rect 119804 141364 119856 141370
rect 119804 141306 119856 141312
rect 119528 140752 119580 140758
rect 119528 140694 119580 140700
rect 119344 140684 119396 140690
rect 119344 140626 119396 140632
rect 119252 140480 119304 140486
rect 119252 140422 119304 140428
rect 119160 140072 119212 140078
rect 119160 140014 119212 140020
rect 119172 80102 119200 140014
rect 119160 80096 119212 80102
rect 119160 80038 119212 80044
rect 119264 79082 119292 140422
rect 119356 79218 119384 140626
rect 119436 140412 119488 140418
rect 119436 140354 119488 140360
rect 119344 79212 119396 79218
rect 119344 79154 119396 79160
rect 119252 79076 119304 79082
rect 119252 79018 119304 79024
rect 119448 76770 119476 140354
rect 119436 76764 119488 76770
rect 119436 76706 119488 76712
rect 119540 75857 119568 140694
rect 119804 139868 119856 139874
rect 119804 139810 119856 139816
rect 119618 138680 119674 138689
rect 119618 138615 119674 138624
rect 119526 75848 119582 75857
rect 119526 75783 119582 75792
rect 119068 71324 119120 71330
rect 119068 71266 119120 71272
rect 119632 70378 119660 138615
rect 119620 70372 119672 70378
rect 119620 70314 119672 70320
rect 119816 69698 119844 139810
rect 120000 73030 120028 200631
rect 120448 148844 120500 148850
rect 120448 148786 120500 148792
rect 120080 78668 120132 78674
rect 120080 78610 120132 78616
rect 120092 75206 120120 78610
rect 120080 75200 120132 75206
rect 120080 75142 120132 75148
rect 119988 73024 120040 73030
rect 119988 72966 120040 72972
rect 120460 70242 120488 148786
rect 120540 144968 120592 144974
rect 120540 144910 120592 144916
rect 120552 97986 120580 144910
rect 120736 142118 120764 259422
rect 120828 142225 120856 260782
rect 120920 143138 120948 263774
rect 121000 263628 121052 263634
rect 121000 263570 121052 263576
rect 120908 143132 120960 143138
rect 120908 143074 120960 143080
rect 121012 142866 121040 263570
rect 132040 263084 132092 263090
rect 132040 263026 132092 263032
rect 127624 262948 127676 262954
rect 127624 262890 127676 262896
rect 131120 262948 131172 262954
rect 131120 262890 131172 262896
rect 131764 262948 131816 262954
rect 131764 262890 131816 262896
rect 125968 262472 126020 262478
rect 125968 262414 126020 262420
rect 122748 262268 122800 262274
rect 122748 262210 122800 262216
rect 122760 260710 122788 262210
rect 125600 260908 125652 260914
rect 125600 260850 125652 260856
rect 123208 260840 123260 260846
rect 123208 260782 123260 260788
rect 122840 260772 122892 260778
rect 122840 260714 122892 260720
rect 122748 260704 122800 260710
rect 122748 260646 122800 260652
rect 122852 259978 122880 260714
rect 123220 259978 123248 260782
rect 124312 260704 124364 260710
rect 124312 260646 124364 260652
rect 123760 260024 123812 260030
rect 122852 259950 123004 259978
rect 123220 259950 123556 259978
rect 124324 259978 124352 260646
rect 125612 259978 125640 260850
rect 125980 259978 126008 262414
rect 127348 261384 127400 261390
rect 127348 261326 127400 261332
rect 127360 261186 127388 261326
rect 127072 261180 127124 261186
rect 127072 261122 127124 261128
rect 127348 261180 127400 261186
rect 127348 261122 127400 261128
rect 127084 259978 127112 261122
rect 127636 259978 127664 262890
rect 131132 262818 131160 262890
rect 131120 262812 131172 262818
rect 131120 262754 131172 262760
rect 131120 262676 131172 262682
rect 131120 262618 131172 262624
rect 129280 262404 129332 262410
rect 129280 262346 129332 262352
rect 128728 261112 128780 261118
rect 128728 261054 128780 261060
rect 128740 259978 128768 261054
rect 129292 259978 129320 262346
rect 129830 262304 129886 262313
rect 129830 262239 129886 262248
rect 129844 261594 129872 262239
rect 129832 261588 129884 261594
rect 129832 261530 129884 261536
rect 129844 259978 129872 261530
rect 131132 261458 131160 262618
rect 131120 261452 131172 261458
rect 131120 261394 131172 261400
rect 130384 261044 130436 261050
rect 130384 260986 130436 260992
rect 130396 259978 130424 260986
rect 131132 259978 131160 261394
rect 131776 259978 131804 262890
rect 132052 261089 132080 263026
rect 132868 261180 132920 261186
rect 132868 261122 132920 261128
rect 132038 261080 132094 261089
rect 132038 261015 132094 261024
rect 132052 259978 132080 261015
rect 123812 259972 124108 259978
rect 123760 259966 124108 259972
rect 123772 259950 124108 259966
rect 124324 259950 124660 259978
rect 125612 259950 125764 259978
rect 125980 259950 126316 259978
rect 127084 259950 127420 259978
rect 127636 259950 127972 259978
rect 128740 259950 129076 259978
rect 129292 259950 129628 259978
rect 129844 259950 130180 259978
rect 130396 259950 130732 259978
rect 131132 259950 131284 259978
rect 131776 259950 131836 259978
rect 132052 259950 132388 259978
rect 128372 259690 128524 259706
rect 128360 259684 128524 259690
rect 128412 259678 128524 259684
rect 128360 259626 128412 259632
rect 132880 259570 132908 261122
rect 133156 259978 133184 263842
rect 134340 261248 134392 261254
rect 134340 261190 134392 261196
rect 134352 260438 134380 261190
rect 134340 260432 134392 260438
rect 134340 260374 134392 260380
rect 134352 259978 134380 260374
rect 133156 259950 133492 259978
rect 134044 259950 134380 259978
rect 134444 259978 134472 263978
rect 134536 262750 134564 324294
rect 134616 298172 134668 298178
rect 134616 298114 134668 298120
rect 134628 264042 134656 298114
rect 134616 264036 134668 264042
rect 134616 263978 134668 263984
rect 134524 262744 134576 262750
rect 134524 262686 134576 262692
rect 134800 262744 134852 262750
rect 134800 262686 134852 262692
rect 134812 259978 134840 262686
rect 135272 260234 135300 351902
rect 135904 311908 135956 311914
rect 135904 311850 135956 311856
rect 135916 265169 135944 311850
rect 137284 286340 137336 286346
rect 137284 286282 137336 286288
rect 137296 267734 137324 286282
rect 137204 267706 137324 267734
rect 135902 265160 135958 265169
rect 135902 265095 135958 265104
rect 135260 260228 135312 260234
rect 135260 260170 135312 260176
rect 134444 259950 134596 259978
rect 134812 259950 135148 259978
rect 135272 259962 135300 260170
rect 135916 259978 135944 265095
rect 137204 263702 137232 267706
rect 137836 267028 137888 267034
rect 137836 266970 137888 266976
rect 137848 264110 137876 266970
rect 137836 264104 137888 264110
rect 137836 264046 137888 264052
rect 137192 263696 137244 263702
rect 137192 263638 137244 263644
rect 136226 260228 136278 260234
rect 136226 260170 136278 260176
rect 135260 259956 135312 259962
rect 135700 259950 135944 259978
rect 136238 259964 136266 260170
rect 137204 259978 137232 263638
rect 137468 263560 137520 263566
rect 137468 263502 137520 263508
rect 137480 260953 137508 263502
rect 137466 260944 137522 260953
rect 137466 260879 137522 260888
rect 136804 259950 137232 259978
rect 135260 259898 135312 259904
rect 137480 259842 137508 260879
rect 137356 259814 137508 259842
rect 137848 259842 137876 264046
rect 138676 262857 138704 430578
rect 138756 418192 138808 418198
rect 138756 418134 138808 418140
rect 138768 265033 138796 418134
rect 139596 267734 139624 484366
rect 140044 470620 140096 470626
rect 140044 470562 140096 470568
rect 140056 267734 140084 470562
rect 140780 280832 140832 280838
rect 140780 280774 140832 280780
rect 139596 267706 139716 267734
rect 140056 267706 140360 267734
rect 138754 265024 138810 265033
rect 138754 264959 138810 264968
rect 138662 262848 138718 262857
rect 138662 262783 138718 262792
rect 138676 259978 138704 262783
rect 138460 259950 138704 259978
rect 138768 259978 138796 264959
rect 139400 264308 139452 264314
rect 139400 264250 139452 264256
rect 139412 263974 139440 264250
rect 139400 263968 139452 263974
rect 139400 263910 139452 263916
rect 139412 259978 139440 263910
rect 139688 260409 139716 267706
rect 140332 262721 140360 267706
rect 140318 262712 140374 262721
rect 140318 262647 140374 262656
rect 139674 260400 139730 260409
rect 139674 260335 139730 260344
rect 139688 259978 139716 260335
rect 140332 259978 140360 262647
rect 140792 260137 140820 280774
rect 141424 265736 141476 265742
rect 141424 265678 141476 265684
rect 141436 263838 141464 265678
rect 141424 263832 141476 263838
rect 141424 263774 141476 263780
rect 140778 260128 140834 260137
rect 140778 260063 140834 260072
rect 141436 259978 141464 263774
rect 142252 262540 142304 262546
rect 142252 262482 142304 262488
rect 141744 260128 141800 260137
rect 141744 260063 141800 260072
rect 138768 259950 139012 259978
rect 139412 259950 139564 259978
rect 139688 259950 140116 259978
rect 140332 259950 140668 259978
rect 141220 259950 141464 259978
rect 141758 259964 141786 260063
rect 142264 259978 142292 262482
rect 142448 260137 142476 590650
rect 142804 563100 142856 563106
rect 142804 563042 142856 563048
rect 142816 267734 142844 563042
rect 142896 524476 142948 524482
rect 142896 524418 142948 524424
rect 142632 267706 142844 267734
rect 142632 263770 142660 267706
rect 142620 263764 142672 263770
rect 142620 263706 142672 263712
rect 142434 260128 142490 260137
rect 142434 260063 142490 260072
rect 142632 259978 142660 263706
rect 142908 262546 142936 524418
rect 142896 262540 142948 262546
rect 142896 262482 142948 262488
rect 143644 260273 143672 616830
rect 144184 576904 144236 576910
rect 144184 576846 144236 576852
rect 144196 262614 144224 576846
rect 145564 289128 145616 289134
rect 145564 289070 145616 289076
rect 144920 282192 144972 282198
rect 144920 282134 144972 282140
rect 144184 262608 144236 262614
rect 144184 262550 144236 262556
rect 143630 260264 143686 260273
rect 143630 260199 143686 260208
rect 143400 260128 143456 260137
rect 143400 260063 143456 260072
rect 142264 259950 142324 259978
rect 142632 259950 142876 259978
rect 143414 259964 143442 260063
rect 144196 259978 144224 262550
rect 144504 260264 144560 260273
rect 144504 260199 144560 260208
rect 143980 259950 144224 259978
rect 144518 259964 144546 260199
rect 144932 259978 144960 282134
rect 145576 263673 145604 289070
rect 146208 268388 146260 268394
rect 146208 268330 146260 268336
rect 146220 263945 146248 268330
rect 146206 263936 146262 263945
rect 146206 263871 146262 263880
rect 145286 263664 145342 263673
rect 145286 263599 145342 263608
rect 145562 263664 145618 263673
rect 145562 263599 145618 263608
rect 145300 259978 145328 263599
rect 146220 260250 146248 263871
rect 146174 260222 146248 260250
rect 144932 259950 145084 259978
rect 145300 259950 145636 259978
rect 146174 259964 146202 260222
rect 146312 259978 146340 696934
rect 146944 683188 146996 683194
rect 146944 683130 146996 683136
rect 146956 262585 146984 683130
rect 147680 282940 147732 282946
rect 147680 282882 147732 282888
rect 147692 263498 147720 282882
rect 147772 269816 147824 269822
rect 147772 269758 147824 269764
rect 147784 263809 147812 269758
rect 148336 267734 148364 700266
rect 149704 345092 149756 345098
rect 149704 345034 149756 345040
rect 149060 287700 149112 287706
rect 149060 287642 149112 287648
rect 148336 267706 148548 267734
rect 147770 263800 147826 263809
rect 147770 263735 147826 263744
rect 147680 263492 147732 263498
rect 147680 263434 147732 263440
rect 146942 262576 146998 262585
rect 146942 262511 146998 262520
rect 146956 259978 146984 262511
rect 147784 259978 147812 263735
rect 148048 263492 148100 263498
rect 148048 263434 148100 263440
rect 148060 259978 148088 263434
rect 148520 262993 148548 267706
rect 148506 262984 148562 262993
rect 148506 262919 148562 262928
rect 148520 259978 148548 262919
rect 146312 259950 146740 259978
rect 146956 259950 147292 259978
rect 147784 259950 147844 259978
rect 148060 259950 148396 259978
rect 148520 259950 148948 259978
rect 144932 259865 144960 259950
rect 144918 259856 144974 259865
rect 137848 259814 137908 259842
rect 144918 259791 144974 259800
rect 146496 259729 146524 259950
rect 146482 259720 146538 259729
rect 146482 259655 146538 259664
rect 149072 259593 149100 287642
rect 149152 271176 149204 271182
rect 149152 271118 149204 271124
rect 149164 259978 149192 271118
rect 149716 264382 149744 345034
rect 150440 284980 150492 284986
rect 150440 284922 150492 284928
rect 149704 264376 149756 264382
rect 149704 264318 149756 264324
rect 149164 259950 149500 259978
rect 149164 259894 149192 259950
rect 149152 259888 149204 259894
rect 149152 259830 149204 259836
rect 150452 259826 150480 284922
rect 151084 275324 151136 275330
rect 151084 275266 151136 275272
rect 151096 263634 151124 275266
rect 151820 273284 151872 273290
rect 151820 273226 151872 273232
rect 151832 267734 151860 273226
rect 151832 267706 152412 267734
rect 152188 264988 152240 264994
rect 152188 264930 152240 264936
rect 151084 263628 151136 263634
rect 151084 263570 151136 263576
rect 150530 262440 150586 262449
rect 150530 262375 150586 262384
rect 150544 259978 150572 262375
rect 151096 259978 151124 263570
rect 152200 259978 152228 264930
rect 152384 259978 152412 267706
rect 152476 264994 152504 700334
rect 152464 264988 152516 264994
rect 152464 264930 152516 264936
rect 153212 262750 153240 702406
rect 157340 700868 157392 700874
rect 157340 700810 157392 700816
rect 155960 700800 156012 700806
rect 155960 700742 156012 700748
rect 154580 700664 154632 700670
rect 154580 700606 154632 700612
rect 153292 700460 153344 700466
rect 153292 700402 153344 700408
rect 153200 262744 153252 262750
rect 153200 262686 153252 262692
rect 153304 259978 153332 700402
rect 153382 276040 153438 276049
rect 153382 275975 153438 275984
rect 153396 267734 153424 275975
rect 153396 267706 154068 267734
rect 153844 262676 153896 262682
rect 153844 262618 153896 262624
rect 153856 259978 153884 262618
rect 154040 259978 154068 267706
rect 154592 259978 154620 700606
rect 155868 262608 155920 262614
rect 155868 262550 155920 262556
rect 155880 259978 155908 262550
rect 155972 260234 156000 700742
rect 156050 277536 156106 277545
rect 156050 277471 156106 277480
rect 155960 260228 156012 260234
rect 155960 260170 156012 260176
rect 150544 259950 150604 259978
rect 151096 259950 151156 259978
rect 152200 259950 152260 259978
rect 152384 259950 152812 259978
rect 153304 259950 153364 259978
rect 153856 259950 153916 259978
rect 154040 259950 154468 259978
rect 154592 259950 155264 259978
rect 155572 259950 155908 259978
rect 156064 259978 156092 277471
rect 157156 262540 157208 262546
rect 157156 262482 157208 262488
rect 156650 260228 156702 260234
rect 156650 260170 156702 260176
rect 156662 259978 156690 260170
rect 157168 259978 157196 262482
rect 157352 260273 157380 700810
rect 160744 700732 160796 700738
rect 160744 700674 160796 700680
rect 157432 450560 157484 450566
rect 157432 450502 157484 450508
rect 157338 260264 157394 260273
rect 157338 260199 157394 260208
rect 157444 259978 157472 450502
rect 160100 279472 160152 279478
rect 160100 279414 160152 279420
rect 158812 269884 158864 269890
rect 158812 269826 158864 269832
rect 158720 264240 158772 264246
rect 158720 264182 158772 264188
rect 158732 263634 158760 264182
rect 158720 263628 158772 263634
rect 158720 263570 158772 263576
rect 158720 262744 158772 262750
rect 158824 262721 158852 269826
rect 159364 263628 159416 263634
rect 159364 263570 159416 263576
rect 158720 262686 158772 262692
rect 158810 262712 158866 262721
rect 158732 261118 158760 262686
rect 158810 262647 158866 262656
rect 158720 261112 158772 261118
rect 158720 261054 158772 261060
rect 158304 260264 158360 260273
rect 158304 260199 158360 260208
rect 156064 259950 156124 259978
rect 156662 259964 157012 259978
rect 156676 259950 157012 259964
rect 157168 259950 157228 259978
rect 157444 259950 158116 259978
rect 153304 259842 153332 259950
rect 151372 259826 151708 259842
rect 150440 259820 150492 259826
rect 150440 259762 150492 259768
rect 151360 259820 151708 259826
rect 151412 259814 151708 259820
rect 153212 259814 153332 259842
rect 151360 259762 151412 259768
rect 153212 259758 153240 259814
rect 153200 259752 153252 259758
rect 153200 259694 153252 259700
rect 155236 259593 155264 259950
rect 156984 259894 157012 259950
rect 156972 259888 157024 259894
rect 156972 259830 157024 259836
rect 158088 259758 158116 259950
rect 158076 259752 158128 259758
rect 158076 259694 158128 259700
rect 158318 259706 158346 260199
rect 158732 259978 158760 261054
rect 159376 259978 159404 263570
rect 159914 262712 159970 262721
rect 159914 262647 159970 262656
rect 159928 259978 159956 262647
rect 160112 260001 160140 279414
rect 160756 267734 160784 700674
rect 162216 700596 162268 700602
rect 162216 700538 162268 700544
rect 162124 700528 162176 700534
rect 162124 700470 162176 700476
rect 161480 683256 161532 683262
rect 161480 683198 161532 683204
rect 160756 267706 160876 267734
rect 160848 264994 160876 267706
rect 160836 264988 160888 264994
rect 160836 264930 160888 264936
rect 160098 259992 160154 260001
rect 158732 259950 158884 259978
rect 159376 259950 159436 259978
rect 159928 259950 159988 259978
rect 160848 259978 160876 264930
rect 161492 260817 161520 683198
rect 162136 267734 162164 700470
rect 162044 267706 162164 267734
rect 162044 262449 162072 267706
rect 162228 265577 162256 700538
rect 163504 670744 163556 670750
rect 163504 670686 163556 670692
rect 162214 265568 162270 265577
rect 162214 265503 162270 265512
rect 162030 262440 162086 262449
rect 162030 262375 162086 262384
rect 161478 260808 161534 260817
rect 161478 260743 161534 260752
rect 160540 259950 160876 259978
rect 160926 259992 160982 260001
rect 160098 259927 160154 259936
rect 162044 259978 162072 262375
rect 162228 260250 162256 265503
rect 163516 265169 163544 670686
rect 163596 656940 163648 656946
rect 163596 656882 163648 656888
rect 163502 265160 163558 265169
rect 163502 265095 163558 265104
rect 163410 263256 163466 263265
rect 163410 263191 163466 263200
rect 163424 262585 163452 263191
rect 163410 262576 163466 262585
rect 163410 262511 163466 262520
rect 162674 260808 162730 260817
rect 162674 260743 162730 260752
rect 160982 259950 161092 259978
rect 161644 259950 162072 259978
rect 162182 260222 162256 260250
rect 162182 259964 162210 260222
rect 160926 259927 160982 259936
rect 162582 259856 162638 259865
rect 162688 259842 162716 260743
rect 163424 259978 163452 262511
rect 163300 259950 163452 259978
rect 163516 259978 163544 265095
rect 163608 263265 163636 656882
rect 164240 632120 164292 632126
rect 164240 632062 164292 632068
rect 163594 263256 163650 263265
rect 163594 263191 163650 263200
rect 164252 259978 164280 632062
rect 164884 618316 164936 618322
rect 164884 618258 164936 618264
rect 164896 265033 164924 618258
rect 164976 605872 165028 605878
rect 164976 605814 165028 605820
rect 164882 265024 164938 265033
rect 164882 264959 164938 264968
rect 164988 262750 165016 605814
rect 165620 579692 165672 579698
rect 165620 579634 165672 579640
rect 165158 265296 165214 265305
rect 165158 265231 165214 265240
rect 165172 265033 165200 265231
rect 165158 265024 165214 265033
rect 165158 264959 165214 264968
rect 164976 262744 165028 262750
rect 164976 262686 165028 262692
rect 164988 260250 165016 262686
rect 164942 260222 165016 260250
rect 164700 260024 164752 260030
rect 163516 259950 163852 259978
rect 164252 259972 164700 259978
rect 164252 259966 164752 259972
rect 164252 259950 164740 259966
rect 164942 259964 164970 260222
rect 165172 259978 165200 264959
rect 165632 259978 165660 579634
rect 167644 565888 167696 565894
rect 167644 565830 167696 565836
rect 166264 553444 166316 553450
rect 166264 553386 166316 553392
rect 166276 262818 166304 553386
rect 167000 527196 167052 527202
rect 167000 527138 167052 527144
rect 166264 262812 166316 262818
rect 166264 262754 166316 262760
rect 166276 259978 166304 262754
rect 167012 260234 167040 527138
rect 167656 267734 167684 565830
rect 167736 501016 167788 501022
rect 167736 500958 167788 500964
rect 167564 267706 167684 267734
rect 167748 267734 167776 500958
rect 169772 450566 169800 702406
rect 202800 700806 202828 703520
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 182824 643136 182876 643142
rect 182824 643078 182876 643084
rect 181444 536852 181496 536858
rect 181444 536794 181496 536800
rect 180064 510672 180116 510678
rect 180064 510614 180116 510620
rect 170404 462392 170456 462398
rect 170404 462334 170456 462340
rect 169760 450560 169812 450566
rect 169760 450502 169812 450508
rect 169760 422340 169812 422346
rect 169760 422282 169812 422288
rect 169024 271244 169076 271250
rect 169024 271186 169076 271192
rect 169036 267734 169064 271186
rect 167748 267706 167868 267734
rect 169036 267706 169156 267734
rect 167458 265568 167514 265577
rect 167458 265503 167514 265512
rect 167472 265169 167500 265503
rect 167564 265441 167592 267706
rect 167550 265432 167606 265441
rect 167550 265367 167606 265376
rect 167458 265160 167514 265169
rect 167458 265095 167514 265104
rect 167000 260228 167052 260234
rect 167000 260170 167052 260176
rect 167564 259978 167592 265367
rect 167840 263022 167868 267706
rect 169128 265130 169156 267706
rect 169208 265668 169260 265674
rect 169208 265610 169260 265616
rect 169116 265124 169168 265130
rect 169116 265066 169168 265072
rect 167828 263016 167880 263022
rect 167828 262958 167880 262964
rect 167690 260228 167742 260234
rect 167690 260170 167742 260176
rect 167702 260098 167730 260170
rect 167690 260092 167742 260098
rect 167690 260034 167742 260040
rect 165172 259950 165508 259978
rect 165632 259962 166212 259978
rect 165632 259956 166224 259962
rect 165632 259950 166172 259956
rect 166276 259950 166612 259978
rect 167164 259950 167592 259978
rect 167702 259964 167730 260034
rect 167840 259978 167868 262958
rect 169128 259978 169156 265066
rect 169220 260166 169248 265610
rect 169772 260234 169800 422282
rect 170220 265328 170272 265334
rect 170220 265270 170272 265276
rect 169760 260228 169812 260234
rect 169760 260170 169812 260176
rect 169208 260160 169260 260166
rect 169208 260102 169260 260108
rect 167840 259950 168268 259978
rect 168820 259950 169156 259978
rect 169220 259978 169248 260102
rect 170232 259978 170260 265270
rect 170416 265062 170444 462334
rect 178684 456816 178736 456822
rect 178684 456758 178736 456764
rect 170496 448588 170548 448594
rect 170496 448530 170548 448536
rect 170508 265334 170536 448530
rect 171784 409896 171836 409902
rect 171784 409838 171836 409844
rect 170496 265328 170548 265334
rect 170496 265270 170548 265276
rect 171692 265260 171744 265266
rect 171692 265202 171744 265208
rect 170404 265056 170456 265062
rect 170404 264998 170456 265004
rect 170680 265056 170732 265062
rect 170680 264998 170732 265004
rect 170692 259978 170720 264998
rect 171002 260228 171054 260234
rect 171002 260170 171054 260176
rect 169220 259950 169372 259978
rect 169924 259950 170260 259978
rect 170476 259950 170720 259978
rect 166172 259898 166224 259904
rect 171014 259842 171042 260170
rect 171704 259978 171732 265202
rect 171796 265198 171824 409838
rect 171876 397520 171928 397526
rect 171876 397462 171928 397468
rect 171888 265538 171916 397462
rect 173900 318844 173952 318850
rect 173900 318786 173952 318792
rect 173164 273964 173216 273970
rect 173164 273906 173216 273912
rect 172520 268456 172572 268462
rect 172520 268398 172572 268404
rect 172532 265606 172560 268398
rect 173176 267734 173204 273906
rect 173176 267706 173388 267734
rect 172520 265600 172572 265606
rect 172520 265542 172572 265548
rect 171876 265532 171928 265538
rect 171876 265474 171928 265480
rect 171888 265266 171916 265474
rect 171876 265260 171928 265266
rect 171876 265202 171928 265208
rect 171784 265192 171836 265198
rect 171784 265134 171836 265140
rect 171580 259950 171732 259978
rect 171796 259978 171824 265134
rect 172532 259978 172560 265542
rect 173360 265266 173388 267706
rect 173348 265260 173400 265266
rect 173348 265202 173400 265208
rect 173164 263696 173216 263702
rect 173164 263638 173216 263644
rect 171796 259950 172132 259978
rect 172532 259950 172684 259978
rect 173176 259842 173204 263638
rect 173360 259978 173388 265202
rect 173440 264376 173492 264382
rect 173440 264318 173492 264324
rect 173452 263702 173480 264318
rect 173440 263696 173492 263702
rect 173440 263638 173492 263644
rect 173912 260506 173940 318786
rect 175924 305040 175976 305046
rect 175924 304982 175976 304988
rect 174544 292596 174596 292602
rect 174544 292538 174596 292544
rect 174556 265470 174584 292538
rect 175936 267734 175964 304982
rect 175844 267706 175964 267734
rect 174544 265464 174596 265470
rect 174544 265406 174596 265412
rect 173900 260500 173952 260506
rect 173900 260442 173952 260448
rect 173912 259978 173940 260442
rect 174556 259978 174584 265406
rect 175844 265402 175872 267706
rect 175924 266416 175976 266422
rect 175924 266358 175976 266364
rect 175832 265396 175884 265402
rect 175832 265338 175884 265344
rect 175844 259978 175872 265338
rect 175936 260302 175964 266358
rect 178696 264314 178724 456758
rect 180076 265742 180104 510614
rect 181456 280838 181484 536794
rect 182836 282198 182864 643078
rect 188344 630692 188396 630698
rect 188344 630634 188396 630640
rect 185584 404388 185636 404394
rect 185584 404330 185636 404336
rect 182824 282192 182876 282198
rect 182824 282134 182876 282140
rect 181444 280832 181496 280838
rect 181444 280774 181496 280780
rect 185596 267034 185624 404330
rect 188356 289134 188384 630634
rect 196624 378208 196676 378214
rect 196624 378150 196676 378156
rect 188344 289128 188396 289134
rect 188344 289070 188396 289076
rect 196636 286346 196664 378150
rect 196624 286340 196676 286346
rect 196624 286282 196676 286288
rect 189448 283620 189500 283626
rect 189448 283562 189500 283568
rect 189460 282946 189488 283562
rect 189080 282940 189132 282946
rect 189080 282882 189132 282888
rect 189448 282940 189500 282946
rect 189448 282882 189500 282888
rect 187700 273964 187752 273970
rect 187700 273906 187752 273912
rect 187712 273290 187740 273906
rect 187700 273284 187752 273290
rect 187700 273226 187752 273232
rect 185584 267028 185636 267034
rect 185584 266970 185636 266976
rect 180064 265736 180116 265742
rect 180064 265678 180116 265684
rect 178684 264308 178736 264314
rect 178684 264250 178736 264256
rect 176752 263152 176804 263158
rect 176752 263094 176804 263100
rect 179236 263152 179288 263158
rect 179236 263094 179288 263100
rect 176200 261316 176252 261322
rect 176200 261258 176252 261264
rect 176212 260982 176240 261258
rect 176764 261186 176792 263094
rect 178408 262880 178460 262886
rect 178408 262822 178460 262828
rect 178420 261526 178448 262822
rect 178408 261520 178460 261526
rect 178408 261462 178460 261468
rect 177304 261316 177356 261322
rect 177304 261258 177356 261264
rect 176752 261180 176804 261186
rect 176752 261122 176804 261128
rect 176200 260976 176252 260982
rect 176200 260918 176252 260924
rect 175924 260296 175976 260302
rect 175924 260238 175976 260244
rect 173360 259950 173788 259978
rect 173912 259950 174340 259978
rect 174556 259950 174892 259978
rect 175444 259950 175872 259978
rect 175936 259978 175964 260238
rect 176212 259978 176240 260918
rect 176764 259978 176792 261122
rect 177316 260370 177344 261258
rect 177304 260364 177356 260370
rect 177304 260306 177356 260312
rect 177316 259978 177344 260306
rect 178420 259978 178448 261462
rect 179248 259978 179276 263094
rect 181812 262472 181864 262478
rect 181812 262414 181864 262420
rect 181260 262336 181312 262342
rect 181260 262278 181312 262284
rect 180524 261248 180576 261254
rect 180524 261190 180576 261196
rect 180536 259978 180564 261190
rect 181272 259978 181300 262278
rect 181824 259978 181852 262414
rect 182916 262404 182968 262410
rect 182916 262346 182968 262352
rect 181996 261044 182048 261050
rect 181996 260986 182048 260992
rect 175936 259950 175996 259978
rect 176212 259950 176548 259978
rect 176764 259950 177100 259978
rect 177316 259950 177652 259978
rect 178420 259950 178756 259978
rect 179248 259950 179308 259978
rect 180412 259950 180564 259978
rect 180964 259950 181300 259978
rect 181516 259950 181852 259978
rect 182008 259978 182036 260986
rect 182928 259978 182956 262346
rect 184572 262268 184624 262274
rect 184572 262210 184624 262216
rect 183468 261384 183520 261390
rect 183468 261326 183520 261332
rect 183480 259978 183508 261326
rect 184020 260908 184072 260914
rect 184020 260850 184072 260856
rect 184032 259978 184060 260850
rect 184584 259978 184612 262210
rect 182008 259950 182068 259978
rect 182620 259950 182956 259978
rect 183172 259950 183508 259978
rect 183724 259950 184060 259978
rect 184276 259950 184612 259978
rect 162638 259814 162748 259842
rect 171014 259828 171180 259842
rect 171028 259826 171180 259828
rect 171028 259820 171192 259826
rect 171028 259814 171140 259820
rect 162582 259791 162638 259800
rect 173176 259814 173236 259842
rect 171140 259762 171192 259768
rect 158626 259720 158682 259729
rect 158318 259692 158626 259706
rect 158332 259678 158626 259692
rect 184828 259690 184980 259706
rect 184828 259684 184992 259690
rect 184828 259678 184940 259684
rect 158626 259655 158682 259664
rect 184940 259626 184992 259632
rect 178040 259616 178092 259622
rect 149058 259584 149114 259593
rect 124876 259542 125212 259570
rect 126532 259554 126868 259570
rect 126520 259548 126868 259554
rect 124876 259486 124904 259542
rect 126572 259542 126868 259548
rect 132880 259542 133276 259570
rect 126520 259490 126572 259496
rect 133248 259486 133276 259542
rect 149058 259519 149114 259528
rect 149794 259584 149850 259593
rect 155222 259584 155278 259593
rect 149850 259542 150052 259570
rect 149794 259519 149850 259528
rect 185674 259584 185730 259593
rect 178092 259564 178204 259570
rect 178040 259558 178204 259564
rect 178052 259542 178204 259558
rect 179860 259554 180196 259570
rect 179860 259548 180208 259554
rect 179860 259542 180156 259548
rect 155222 259519 155278 259528
rect 185380 259542 185674 259570
rect 185674 259519 185730 259528
rect 180156 259490 180208 259496
rect 124864 259480 124916 259486
rect 124864 259422 124916 259428
rect 133236 259480 133288 259486
rect 133236 259422 133288 259428
rect 128912 200728 128964 200734
rect 128912 200670 128964 200676
rect 129280 200728 129332 200734
rect 129280 200670 129332 200676
rect 131580 200728 131632 200734
rect 131580 200670 131632 200676
rect 131672 200728 131724 200734
rect 178776 200728 178828 200734
rect 131672 200670 131724 200676
rect 132038 200696 132094 200705
rect 128084 200592 128136 200598
rect 128084 200534 128136 200540
rect 123944 200388 123996 200394
rect 123944 200330 123996 200336
rect 121092 200320 121144 200326
rect 121092 200262 121144 200268
rect 121000 142860 121052 142866
rect 121000 142802 121052 142808
rect 120814 142216 120870 142225
rect 120814 142151 120870 142160
rect 120724 142112 120776 142118
rect 120724 142054 120776 142060
rect 120816 141568 120868 141574
rect 120816 141510 120868 141516
rect 120632 140004 120684 140010
rect 120632 139946 120684 139952
rect 120540 97980 120592 97986
rect 120540 97922 120592 97928
rect 120644 79150 120672 139946
rect 120724 80912 120776 80918
rect 120724 80854 120776 80860
rect 120736 80714 120764 80854
rect 120724 80708 120776 80714
rect 120724 80650 120776 80656
rect 120632 79144 120684 79150
rect 120632 79086 120684 79092
rect 120828 71398 120856 141510
rect 120908 141500 120960 141506
rect 120908 141442 120960 141448
rect 120816 71392 120868 71398
rect 120816 71334 120868 71340
rect 120448 70236 120500 70242
rect 120448 70178 120500 70184
rect 120920 70174 120948 141442
rect 121000 140548 121052 140554
rect 121000 140490 121052 140496
rect 121012 71262 121040 140490
rect 121104 76809 121132 200262
rect 122748 199368 122800 199374
rect 122748 199310 122800 199316
rect 123850 199336 123906 199345
rect 122564 199300 122616 199306
rect 122564 199242 122616 199248
rect 122472 199232 122524 199238
rect 122472 199174 122524 199180
rect 122380 199164 122432 199170
rect 122380 199106 122432 199112
rect 121184 199096 121236 199102
rect 121184 199038 121236 199044
rect 121090 76800 121146 76809
rect 121090 76735 121146 76744
rect 121196 75449 121224 199038
rect 121276 199028 121328 199034
rect 121276 198970 121328 198976
rect 121288 75546 121316 198970
rect 122104 198280 122156 198286
rect 122104 198222 122156 198228
rect 121368 195288 121420 195294
rect 121368 195230 121420 195236
rect 121380 78674 121408 195230
rect 121920 195016 121972 195022
rect 121920 194958 121972 194964
rect 121736 148300 121788 148306
rect 121736 148242 121788 148248
rect 121748 142202 121776 148242
rect 121932 147801 121960 194958
rect 122012 148708 122064 148714
rect 122012 148650 122064 148656
rect 121918 147792 121974 147801
rect 121918 147727 121974 147736
rect 121748 142174 121960 142202
rect 121932 138014 121960 142174
rect 121748 137986 121960 138014
rect 121642 85232 121698 85241
rect 121642 85167 121698 85176
rect 121656 81054 121684 85167
rect 121644 81048 121696 81054
rect 121644 80990 121696 80996
rect 121368 78668 121420 78674
rect 121368 78610 121420 78616
rect 121276 75540 121328 75546
rect 121276 75482 121328 75488
rect 121182 75440 121238 75449
rect 121182 75375 121238 75384
rect 121000 71256 121052 71262
rect 121000 71198 121052 71204
rect 121748 70310 121776 137986
rect 122024 133362 122052 148650
rect 121840 133334 122052 133362
rect 121840 122834 121868 133334
rect 122116 133226 122144 198222
rect 122196 195220 122248 195226
rect 122196 195162 122248 195168
rect 122024 133198 122144 133226
rect 122024 122890 122052 133198
rect 122208 133090 122236 195162
rect 122288 195152 122340 195158
rect 122288 195094 122340 195100
rect 122116 133062 122236 133090
rect 122116 123026 122144 133062
rect 122194 128480 122250 128489
rect 122194 128415 122250 128424
rect 122208 123185 122236 128415
rect 122194 123176 122250 123185
rect 122194 123111 122250 123120
rect 122116 122998 122236 123026
rect 122024 122862 122144 122890
rect 121840 122806 122052 122834
rect 121918 122768 121974 122777
rect 121918 122703 121974 122712
rect 121932 113393 121960 122703
rect 121918 113384 121974 113393
rect 121918 113319 121974 113328
rect 122024 113174 122052 122806
rect 122116 122777 122144 122862
rect 122102 122768 122158 122777
rect 122102 122703 122158 122712
rect 122208 122618 122236 122998
rect 122116 122590 122236 122618
rect 122116 113370 122144 122590
rect 122194 122496 122250 122505
rect 122194 122431 122250 122440
rect 122208 113529 122236 122431
rect 122194 113520 122250 113529
rect 122194 113455 122250 113464
rect 122116 113342 122236 113370
rect 122102 113248 122158 113257
rect 122102 113183 122158 113192
rect 121840 113146 122052 113174
rect 121840 103514 121868 113146
rect 122116 113098 122144 113183
rect 121932 113070 122144 113098
rect 121932 103578 121960 113070
rect 122208 112962 122236 113342
rect 122116 112934 122236 112962
rect 122116 103714 122144 112934
rect 122194 112840 122250 112849
rect 122194 112775 122250 112784
rect 122208 103873 122236 112775
rect 122194 103864 122250 103873
rect 122194 103799 122250 103808
rect 122116 103686 122236 103714
rect 121932 103550 122144 103578
rect 121840 103486 122052 103514
rect 121918 103320 121974 103329
rect 121918 103255 121974 103264
rect 121932 94081 121960 103255
rect 121918 94072 121974 94081
rect 121918 94007 121974 94016
rect 122024 93854 122052 103486
rect 122116 103465 122144 103550
rect 122102 103456 122158 103465
rect 122102 103391 122158 103400
rect 122208 103306 122236 103686
rect 122116 103278 122236 103306
rect 122116 94058 122144 103278
rect 122194 103184 122250 103193
rect 122194 103119 122250 103128
rect 122208 94217 122236 103119
rect 122194 94208 122250 94217
rect 122194 94143 122250 94152
rect 122116 94030 122236 94058
rect 122102 93936 122158 93945
rect 122102 93871 122158 93880
rect 121840 93826 122052 93854
rect 121840 84810 121868 93826
rect 122116 93786 122144 93871
rect 122024 93758 122144 93786
rect 122024 85241 122052 93758
rect 122208 93650 122236 94030
rect 122116 93622 122236 93650
rect 122010 85232 122066 85241
rect 122010 85167 122066 85176
rect 121840 84782 122052 84810
rect 121920 81252 121972 81258
rect 121920 81194 121972 81200
rect 121932 75177 121960 81194
rect 121918 75168 121974 75177
rect 121918 75103 121974 75112
rect 121736 70304 121788 70310
rect 121736 70246 121788 70252
rect 120908 70168 120960 70174
rect 120908 70110 120960 70116
rect 122024 70106 122052 84782
rect 122116 80054 122144 93622
rect 122194 93528 122250 93537
rect 122194 93463 122250 93472
rect 122208 89729 122236 93463
rect 122194 89720 122250 89729
rect 122194 89655 122250 89664
rect 122300 85082 122328 195094
rect 122392 85105 122420 199106
rect 122208 85054 122328 85082
rect 122378 85096 122434 85105
rect 122208 81258 122236 85054
rect 122378 85031 122434 85040
rect 122484 84946 122512 199174
rect 122300 84918 122512 84946
rect 122196 81252 122248 81258
rect 122196 81194 122248 81200
rect 122116 80026 122236 80054
rect 122208 78334 122236 80026
rect 122196 78328 122248 78334
rect 122196 78270 122248 78276
rect 122300 75206 122328 84918
rect 122378 84688 122434 84697
rect 122378 84623 122434 84632
rect 122392 77178 122420 84623
rect 122470 80336 122526 80345
rect 122470 80271 122526 80280
rect 122380 77172 122432 77178
rect 122380 77114 122432 77120
rect 122288 75200 122340 75206
rect 122288 75142 122340 75148
rect 122484 74633 122512 80271
rect 122576 75478 122604 199242
rect 122656 198756 122708 198762
rect 122656 198698 122708 198704
rect 122564 75472 122616 75478
rect 122564 75414 122616 75420
rect 122668 75313 122696 198698
rect 122654 75304 122710 75313
rect 122654 75239 122710 75248
rect 122470 74624 122526 74633
rect 122470 74559 122526 74568
rect 122760 72418 122788 199310
rect 123850 199271 123906 199280
rect 123758 199200 123814 199209
rect 123758 199135 123814 199144
rect 123116 198620 123168 198626
rect 123116 198562 123168 198568
rect 123024 196512 123076 196518
rect 123024 196454 123076 196460
rect 122840 79620 122892 79626
rect 122840 79562 122892 79568
rect 122748 72412 122800 72418
rect 122748 72354 122800 72360
rect 122852 71738 122880 79562
rect 123036 78130 123064 196454
rect 123128 81122 123156 198562
rect 123668 197668 123720 197674
rect 123668 197610 123720 197616
rect 123392 193656 123444 193662
rect 123392 193598 123444 193604
rect 123206 139632 123262 139641
rect 123206 139567 123262 139576
rect 123116 81116 123168 81122
rect 123116 81058 123168 81064
rect 123024 78124 123076 78130
rect 123024 78066 123076 78072
rect 123220 74050 123248 139567
rect 123298 138816 123354 138825
rect 123298 138751 123354 138760
rect 123208 74044 123260 74050
rect 123208 73986 123260 73992
rect 123312 71738 123340 138751
rect 123404 78266 123432 193598
rect 123484 141364 123536 141370
rect 123484 141306 123536 141312
rect 123496 140321 123524 141306
rect 123482 140312 123538 140321
rect 123482 140247 123538 140256
rect 123496 139890 123524 140247
rect 123496 139862 123556 139890
rect 123680 79286 123708 197610
rect 123668 79280 123720 79286
rect 123668 79222 123720 79228
rect 123392 78260 123444 78266
rect 123392 78202 123444 78208
rect 123772 73098 123800 199135
rect 123760 73092 123812 73098
rect 123760 73034 123812 73040
rect 123864 72593 123892 199271
rect 123850 72584 123906 72593
rect 123956 72554 123984 200330
rect 127622 200288 127678 200297
rect 127622 200223 127678 200232
rect 126152 199708 126204 199714
rect 126152 199650 126204 199656
rect 126164 198014 126192 199650
rect 126336 198824 126388 198830
rect 126336 198766 126388 198772
rect 126152 198008 126204 198014
rect 126152 197950 126204 197956
rect 124864 196580 124916 196586
rect 124864 196522 124916 196528
rect 124312 142724 124364 142730
rect 124312 142666 124364 142672
rect 124034 142216 124090 142225
rect 124034 142151 124090 142160
rect 124048 139890 124076 142151
rect 124048 139862 124108 139890
rect 124324 139482 124352 142666
rect 124772 140684 124824 140690
rect 124772 140626 124824 140632
rect 124784 139942 124812 140626
rect 124772 139936 124824 139942
rect 124772 139878 124824 139884
rect 124876 139738 124904 196522
rect 125048 148912 125100 148918
rect 125048 148854 125100 148860
rect 124954 148472 125010 148481
rect 124954 148407 125010 148416
rect 124864 139732 124916 139738
rect 124864 139674 124916 139680
rect 124324 139466 124904 139482
rect 124324 139460 124916 139466
rect 124324 139454 124864 139460
rect 124864 139402 124916 139408
rect 124968 139369 124996 148407
rect 125060 139641 125088 148854
rect 126348 142154 126376 198766
rect 126796 197804 126848 197810
rect 126796 197746 126848 197752
rect 126704 197736 126756 197742
rect 126704 197678 126756 197684
rect 126716 197441 126744 197678
rect 126702 197432 126758 197441
rect 126702 197367 126758 197376
rect 126428 195084 126480 195090
rect 126428 195026 126480 195032
rect 126164 142126 126376 142154
rect 126060 142112 126112 142118
rect 126060 142054 126112 142060
rect 125508 141296 125560 141302
rect 125508 141238 125560 141244
rect 125520 140865 125548 141238
rect 126072 141166 126100 142054
rect 126060 141160 126112 141166
rect 126060 141102 126112 141108
rect 125506 140856 125562 140865
rect 125506 140791 125562 140800
rect 125520 139890 125548 140791
rect 126072 139890 126100 141102
rect 126164 140078 126192 142126
rect 126244 141772 126296 141778
rect 126244 141714 126296 141720
rect 126256 141001 126284 141714
rect 126242 140992 126298 141001
rect 126242 140927 126298 140936
rect 126152 140072 126204 140078
rect 126152 140014 126204 140020
rect 125212 139862 125548 139890
rect 125764 139862 126100 139890
rect 126256 139890 126284 140927
rect 126256 139862 126316 139890
rect 125046 139632 125102 139641
rect 125046 139567 125102 139576
rect 126440 139398 126468 195026
rect 126612 183524 126664 183530
rect 126612 183466 126664 183472
rect 126624 142154 126652 183466
rect 126808 180794 126836 197746
rect 126532 142126 126652 142154
rect 126716 180766 126836 180794
rect 126532 139874 126560 142126
rect 126610 140312 126666 140321
rect 126610 140247 126666 140256
rect 126624 140078 126652 140247
rect 126612 140072 126664 140078
rect 126612 140014 126664 140020
rect 126520 139868 126572 139874
rect 126520 139810 126572 139816
rect 126152 139392 126204 139398
rect 124954 139360 125010 139369
rect 124954 139295 125010 139304
rect 126150 139360 126152 139369
rect 126428 139392 126480 139398
rect 126204 139360 126206 139369
rect 126716 139369 126744 180766
rect 127532 147280 127584 147286
rect 127532 147222 127584 147228
rect 127544 146334 127572 147222
rect 127532 146328 127584 146334
rect 127532 146270 127584 146276
rect 126796 141976 126848 141982
rect 126796 141918 126848 141924
rect 126808 140894 126836 141918
rect 127348 141840 127400 141846
rect 127348 141782 127400 141788
rect 126796 140888 126848 140894
rect 126796 140830 126848 140836
rect 126808 139890 126836 140830
rect 127360 139890 127388 141782
rect 127544 139890 127572 146270
rect 127636 140185 127664 200223
rect 128096 193905 128124 200534
rect 128360 199912 128412 199918
rect 128360 199854 128412 199860
rect 128268 197940 128320 197946
rect 128268 197882 128320 197888
rect 128082 193896 128138 193905
rect 128082 193831 128138 193840
rect 127716 193180 127768 193186
rect 127716 193122 127768 193128
rect 127728 143478 127756 193122
rect 127808 192364 127860 192370
rect 127808 192306 127860 192312
rect 127820 146266 127848 192306
rect 127808 146260 127860 146266
rect 127808 146202 127860 146208
rect 127716 143472 127768 143478
rect 127716 143414 127768 143420
rect 127622 140176 127678 140185
rect 127622 140111 127678 140120
rect 126808 139862 126868 139890
rect 127360 139876 127420 139890
rect 127360 139862 127434 139876
rect 127544 139862 127972 139890
rect 127406 139754 127434 139862
rect 127406 139740 127572 139754
rect 127420 139726 127572 139740
rect 127544 139534 127572 139726
rect 127532 139528 127584 139534
rect 127532 139470 127584 139476
rect 128280 139369 128308 197882
rect 128372 193730 128400 199854
rect 128544 199844 128596 199850
rect 128544 199786 128596 199792
rect 128556 198422 128584 199786
rect 128544 198416 128596 198422
rect 128544 198358 128596 198364
rect 128924 198082 128952 200670
rect 129096 199980 129148 199986
rect 129096 199922 129148 199928
rect 129002 199880 129058 199889
rect 129002 199815 129058 199824
rect 129016 198558 129044 199815
rect 129004 198552 129056 198558
rect 129004 198494 129056 198500
rect 128912 198076 128964 198082
rect 128912 198018 128964 198024
rect 129002 196480 129058 196489
rect 129002 196415 129058 196424
rect 128728 196036 128780 196042
rect 128728 195978 128780 195984
rect 128740 195401 128768 195978
rect 128726 195392 128782 195401
rect 128726 195327 128782 195336
rect 128360 193724 128412 193730
rect 128360 193666 128412 193672
rect 128360 147144 128412 147150
rect 128360 147086 128412 147092
rect 128372 146402 128400 147086
rect 128360 146396 128412 146402
rect 128360 146338 128412 146344
rect 128372 140758 128400 146338
rect 128912 146192 128964 146198
rect 128912 146134 128964 146140
rect 128924 143546 128952 146134
rect 128452 143540 128504 143546
rect 128452 143482 128504 143488
rect 128912 143540 128964 143546
rect 128912 143482 128964 143488
rect 128360 140752 128412 140758
rect 128360 140694 128412 140700
rect 128464 139618 128492 143482
rect 128924 139890 128952 143482
rect 129016 140690 129044 196415
rect 129004 140684 129056 140690
rect 129004 140626 129056 140632
rect 129108 140622 129136 199922
rect 129292 199073 129320 200670
rect 130476 200456 130528 200462
rect 130474 200424 130476 200433
rect 130528 200424 130530 200433
rect 130474 200359 130530 200368
rect 131302 200424 131358 200433
rect 131302 200359 131358 200368
rect 131316 200161 131344 200359
rect 131488 200252 131540 200258
rect 131488 200194 131540 200200
rect 130014 200152 130070 200161
rect 130014 200087 130070 200096
rect 131302 200152 131358 200161
rect 131302 200087 131358 200096
rect 129554 199608 129610 199617
rect 129554 199543 129610 199552
rect 129278 199064 129334 199073
rect 129278 198999 129334 199008
rect 129568 198966 129596 199543
rect 130028 199374 130056 200087
rect 131500 199578 131528 200194
rect 131592 199753 131620 200670
rect 131684 200161 131712 200670
rect 132038 200631 132094 200640
rect 132222 200696 132278 200705
rect 132222 200631 132224 200640
rect 132052 200598 132080 200631
rect 132276 200631 132278 200640
rect 178682 200696 178738 200705
rect 178776 200670 178828 200676
rect 178682 200631 178738 200640
rect 132224 200602 132276 200608
rect 131948 200592 132000 200598
rect 131948 200534 132000 200540
rect 132040 200592 132092 200598
rect 132040 200534 132092 200540
rect 131764 200524 131816 200530
rect 131764 200466 131816 200472
rect 131776 200190 131804 200466
rect 131856 200456 131908 200462
rect 131856 200398 131908 200404
rect 131764 200184 131816 200190
rect 131670 200152 131726 200161
rect 131764 200126 131816 200132
rect 131868 200122 131896 200398
rect 131670 200087 131726 200096
rect 131856 200116 131908 200122
rect 131856 200058 131908 200064
rect 131762 199880 131818 199889
rect 131762 199815 131818 199824
rect 131776 199782 131804 199815
rect 131764 199776 131816 199782
rect 131578 199744 131634 199753
rect 131764 199718 131816 199724
rect 131578 199679 131634 199688
rect 131960 199646 131988 200534
rect 178314 200152 178370 200161
rect 132052 200110 132388 200138
rect 131856 199640 131908 199646
rect 131856 199582 131908 199588
rect 131948 199640 132000 199646
rect 131948 199582 132000 199588
rect 131488 199572 131540 199578
rect 131488 199514 131540 199520
rect 130016 199368 130068 199374
rect 130016 199310 130068 199316
rect 129556 198960 129608 198966
rect 129556 198902 129608 198908
rect 129188 198892 129240 198898
rect 129188 198834 129240 198840
rect 129096 140616 129148 140622
rect 129096 140558 129148 140564
rect 129200 140010 129228 198834
rect 131764 198552 131816 198558
rect 131764 198494 131816 198500
rect 130384 198416 130436 198422
rect 130384 198358 130436 198364
rect 129280 196444 129332 196450
rect 129280 196386 129332 196392
rect 129292 151814 129320 196386
rect 129292 151786 129596 151814
rect 129464 141160 129516 141166
rect 129464 141102 129516 141108
rect 129476 140894 129504 141102
rect 129464 140888 129516 140894
rect 129464 140830 129516 140836
rect 129280 140752 129332 140758
rect 129280 140694 129332 140700
rect 129188 140004 129240 140010
rect 129188 139946 129240 139952
rect 129292 139890 129320 140694
rect 129568 140162 129596 151786
rect 130290 146296 130346 146305
rect 130290 146231 130346 146240
rect 129830 146160 129886 146169
rect 129830 146095 129886 146104
rect 129924 146124 129976 146130
rect 129738 146024 129794 146033
rect 129738 145959 129794 145968
rect 129752 143478 129780 145959
rect 129740 143472 129792 143478
rect 129740 143414 129792 143420
rect 129844 142798 129872 146095
rect 129924 146066 129976 146072
rect 129832 142792 129884 142798
rect 129832 142734 129884 142740
rect 129936 142254 129964 146066
rect 130200 144220 130252 144226
rect 130200 144162 130252 144168
rect 129924 142248 129976 142254
rect 129924 142190 129976 142196
rect 130212 140162 130240 144162
rect 129476 140134 129596 140162
rect 130166 140134 130240 140162
rect 129476 140010 129504 140134
rect 129464 140004 129516 140010
rect 129464 139946 129516 139952
rect 128924 139862 129076 139890
rect 129292 139862 129628 139890
rect 130166 139876 130194 140134
rect 130304 139890 130332 146231
rect 130396 144770 130424 198358
rect 130474 197160 130530 197169
rect 130474 197095 130530 197104
rect 130384 144764 130436 144770
rect 130384 144706 130436 144712
rect 130488 142730 130516 197095
rect 130568 192296 130620 192302
rect 130568 192238 130620 192244
rect 130580 144702 130608 192238
rect 131304 146056 131356 146062
rect 131304 145998 131356 146004
rect 130568 144696 130620 144702
rect 130568 144638 130620 144644
rect 131212 144288 131264 144294
rect 131212 144230 131264 144236
rect 130476 142724 130528 142730
rect 130476 142666 130528 142672
rect 131224 139890 131252 144230
rect 131316 140758 131344 145998
rect 131580 145988 131632 145994
rect 131580 145930 131632 145936
rect 131592 143342 131620 145930
rect 131776 145926 131804 198494
rect 131868 198490 131896 199582
rect 131856 198484 131908 198490
rect 131856 198426 131908 198432
rect 131856 195356 131908 195362
rect 131856 195298 131908 195304
rect 131868 147218 131896 195298
rect 132052 195294 132080 200110
rect 132222 200016 132278 200025
rect 132222 199951 132224 199960
rect 132276 199951 132278 199960
rect 132224 199922 132276 199928
rect 132130 199880 132186 199889
rect 132466 199832 132494 200124
rect 132558 199918 132586 200124
rect 132650 199918 132678 200124
rect 132546 199912 132598 199918
rect 132546 199854 132598 199860
rect 132638 199912 132690 199918
rect 132638 199854 132690 199860
rect 132130 199815 132132 199824
rect 132184 199815 132186 199824
rect 132132 199786 132184 199792
rect 132420 199804 132494 199832
rect 132224 197872 132276 197878
rect 132224 197814 132276 197820
rect 132040 195288 132092 195294
rect 132040 195230 132092 195236
rect 131856 147212 131908 147218
rect 131856 147154 131908 147160
rect 131764 145920 131816 145926
rect 131764 145862 131816 145868
rect 131488 143336 131540 143342
rect 131488 143278 131540 143284
rect 131580 143336 131632 143342
rect 131580 143278 131632 143284
rect 131304 140752 131356 140758
rect 131304 140694 131356 140700
rect 131500 139890 131528 143278
rect 130304 139862 130732 139890
rect 131224 139862 131284 139890
rect 131500 139862 131836 139890
rect 128464 139602 128860 139618
rect 128464 139596 128872 139602
rect 128464 139590 128820 139596
rect 128820 139538 128872 139544
rect 132236 139369 132264 197814
rect 132420 196081 132448 199804
rect 132742 199628 132770 200124
rect 132834 199730 132862 200124
rect 132926 199889 132954 200124
rect 133018 199918 133046 200124
rect 133006 199912 133058 199918
rect 132912 199880 132968 199889
rect 133006 199854 133058 199860
rect 132912 199815 132968 199824
rect 133110 199730 133138 200124
rect 133202 199918 133230 200124
rect 133190 199912 133242 199918
rect 133190 199854 133242 199860
rect 132834 199702 132908 199730
rect 132498 199608 132554 199617
rect 132498 199543 132554 199552
rect 132696 199600 132770 199628
rect 132512 199442 132540 199543
rect 132500 199436 132552 199442
rect 132500 199378 132552 199384
rect 132696 196217 132724 199600
rect 132776 199096 132828 199102
rect 132776 199038 132828 199044
rect 132788 198082 132816 199038
rect 132776 198076 132828 198082
rect 132776 198018 132828 198024
rect 132776 197600 132828 197606
rect 132776 197542 132828 197548
rect 132788 197130 132816 197542
rect 132776 197124 132828 197130
rect 132776 197066 132828 197072
rect 132682 196208 132738 196217
rect 132682 196143 132738 196152
rect 132880 196081 132908 199702
rect 133064 199702 133138 199730
rect 133294 199730 133322 200124
rect 133386 199889 133414 200124
rect 133372 199880 133428 199889
rect 133372 199815 133428 199824
rect 133478 199764 133506 200124
rect 133432 199736 133506 199764
rect 133294 199702 133368 199730
rect 132960 199504 133012 199510
rect 132960 199446 133012 199452
rect 132972 199102 133000 199446
rect 132960 199096 133012 199102
rect 132960 199038 133012 199044
rect 132960 197192 133012 197198
rect 132960 197134 133012 197140
rect 132972 196314 133000 197134
rect 132960 196308 133012 196314
rect 132960 196250 133012 196256
rect 132406 196072 132462 196081
rect 132406 196007 132462 196016
rect 132866 196072 132922 196081
rect 132866 196007 132922 196016
rect 133064 191834 133092 199702
rect 133144 199640 133196 199646
rect 133144 199582 133196 199588
rect 133156 199374 133184 199582
rect 133340 199458 133368 199702
rect 133248 199430 133368 199458
rect 133144 199368 133196 199374
rect 133144 199310 133196 199316
rect 133248 198218 133276 199430
rect 133328 199368 133380 199374
rect 133328 199310 133380 199316
rect 133236 198212 133288 198218
rect 133236 198154 133288 198160
rect 133340 197849 133368 199310
rect 133326 197840 133382 197849
rect 133326 197775 133382 197784
rect 133326 197704 133382 197713
rect 133326 197639 133382 197648
rect 133236 197056 133288 197062
rect 133236 196998 133288 197004
rect 133144 196716 133196 196722
rect 133144 196658 133196 196664
rect 133156 196382 133184 196658
rect 133248 196654 133276 196998
rect 133236 196648 133288 196654
rect 133236 196590 133288 196596
rect 133144 196376 133196 196382
rect 133144 196318 133196 196324
rect 133340 195702 133368 197639
rect 133328 195696 133380 195702
rect 133328 195638 133380 195644
rect 132696 191806 133092 191834
rect 132696 148345 132724 191806
rect 133432 180794 133460 199736
rect 133570 199696 133598 200124
rect 133662 199889 133690 200124
rect 133754 199918 133782 200124
rect 133742 199912 133794 199918
rect 133648 199880 133704 199889
rect 133742 199854 133794 199860
rect 133648 199815 133704 199824
rect 133696 199776 133748 199782
rect 133846 199730 133874 200124
rect 133938 199889 133966 200124
rect 134030 199918 134058 200124
rect 134018 199912 134070 199918
rect 133924 199880 133980 199889
rect 134018 199854 134070 199860
rect 133924 199815 133980 199824
rect 133696 199718 133748 199724
rect 133524 199668 133598 199696
rect 133524 198665 133552 199668
rect 133510 198656 133566 198665
rect 133510 198591 133566 198600
rect 133708 197985 133736 199718
rect 133800 199702 133874 199730
rect 133972 199776 134024 199782
rect 134122 199730 134150 200124
rect 133972 199718 134024 199724
rect 133694 197976 133750 197985
rect 133694 197911 133750 197920
rect 133800 180794 133828 199702
rect 133880 199504 133932 199510
rect 133880 199446 133932 199452
rect 133892 197849 133920 199446
rect 133984 198150 134012 199718
rect 134076 199702 134150 199730
rect 134076 198734 134104 199702
rect 134214 199628 134242 200124
rect 134306 199730 134334 200124
rect 134398 199918 134426 200124
rect 134386 199912 134438 199918
rect 134386 199854 134438 199860
rect 134490 199764 134518 200124
rect 134582 199918 134610 200124
rect 134570 199912 134622 199918
rect 134570 199854 134622 199860
rect 134444 199753 134518 199764
rect 134430 199744 134518 199753
rect 134306 199702 134380 199730
rect 134214 199600 134288 199628
rect 134076 198706 134196 198734
rect 133972 198144 134024 198150
rect 133972 198086 134024 198092
rect 133878 197840 133934 197849
rect 133878 197775 133934 197784
rect 133972 195696 134024 195702
rect 133972 195638 134024 195644
rect 133984 195362 134012 195638
rect 134168 195498 134196 198706
rect 134260 195974 134288 199600
rect 134352 199510 134380 199702
rect 134486 199736 134518 199744
rect 134674 199730 134702 200124
rect 134430 199679 134486 199688
rect 134628 199702 134702 199730
rect 134432 199640 134484 199646
rect 134432 199582 134484 199588
rect 134340 199504 134392 199510
rect 134340 199446 134392 199452
rect 134444 197985 134472 199582
rect 134628 199560 134656 199702
rect 134766 199628 134794 200124
rect 134858 199850 134886 200124
rect 134846 199844 134898 199850
rect 134846 199786 134898 199792
rect 134950 199730 134978 200124
rect 135042 199918 135070 200124
rect 135030 199912 135082 199918
rect 135030 199854 135082 199860
rect 134536 199532 134656 199560
rect 134720 199600 134794 199628
rect 134904 199702 134978 199730
rect 134430 197976 134486 197985
rect 134430 197911 134486 197920
rect 134536 197033 134564 199532
rect 134616 199368 134668 199374
rect 134616 199310 134668 199316
rect 134522 197024 134578 197033
rect 134522 196959 134578 196968
rect 134260 195946 134380 195974
rect 134156 195492 134208 195498
rect 134156 195434 134208 195440
rect 133972 195356 134024 195362
rect 133972 195298 134024 195304
rect 134064 195356 134116 195362
rect 134064 195298 134116 195304
rect 134076 190058 134104 195298
rect 134248 195288 134300 195294
rect 134248 195230 134300 195236
rect 134064 190052 134116 190058
rect 134064 189994 134116 190000
rect 133064 180766 133460 180794
rect 133708 180766 133828 180794
rect 132682 148336 132738 148345
rect 132682 148271 132738 148280
rect 132590 143304 132646 143313
rect 132590 143239 132646 143248
rect 132316 140752 132368 140758
rect 132316 140694 132368 140700
rect 132328 139890 132356 140694
rect 132604 139890 132632 143239
rect 132328 139862 132388 139890
rect 132604 139862 132940 139890
rect 133064 139369 133092 180766
rect 133708 148646 133736 180766
rect 133696 148640 133748 148646
rect 133696 148582 133748 148588
rect 134260 148578 134288 195230
rect 134352 190454 134380 195946
rect 134628 195294 134656 199310
rect 134616 195288 134668 195294
rect 134616 195230 134668 195236
rect 134720 192982 134748 199600
rect 134800 199504 134852 199510
rect 134800 199446 134852 199452
rect 134812 197538 134840 199446
rect 134800 197532 134852 197538
rect 134800 197474 134852 197480
rect 134904 194138 134932 199702
rect 134984 199640 135036 199646
rect 135134 199628 135162 200124
rect 135226 199730 135254 200124
rect 135318 199850 135346 200124
rect 135410 199918 135438 200124
rect 135398 199912 135450 199918
rect 135502 199889 135530 200124
rect 135594 199918 135622 200124
rect 135686 199918 135714 200124
rect 135778 199918 135806 200124
rect 135582 199912 135634 199918
rect 135398 199854 135450 199860
rect 135488 199880 135544 199889
rect 135306 199844 135358 199850
rect 135582 199854 135634 199860
rect 135674 199912 135726 199918
rect 135674 199854 135726 199860
rect 135766 199912 135818 199918
rect 135766 199854 135818 199860
rect 135488 199815 135544 199824
rect 135306 199786 135358 199792
rect 135720 199776 135772 199782
rect 135442 199744 135498 199753
rect 135226 199702 135300 199730
rect 135134 199600 135208 199628
rect 134984 199582 135036 199588
rect 134996 195362 135024 199582
rect 135076 198688 135128 198694
rect 135076 198630 135128 198636
rect 135088 195974 135116 198630
rect 135180 197985 135208 199600
rect 135272 198694 135300 199702
rect 135870 199764 135898 200124
rect 135720 199718 135772 199724
rect 135824 199736 135898 199764
rect 135442 199679 135498 199688
rect 135628 199708 135680 199714
rect 135260 198688 135312 198694
rect 135260 198630 135312 198636
rect 135258 198520 135314 198529
rect 135258 198455 135314 198464
rect 135166 197976 135222 197985
rect 135166 197911 135222 197920
rect 135272 197441 135300 198455
rect 135352 197532 135404 197538
rect 135352 197474 135404 197480
rect 135258 197432 135314 197441
rect 135258 197367 135314 197376
rect 135088 195946 135208 195974
rect 134984 195356 135036 195362
rect 134984 195298 135036 195304
rect 135180 194410 135208 195946
rect 135168 194404 135220 194410
rect 135168 194346 135220 194352
rect 134892 194132 134944 194138
rect 134892 194074 134944 194080
rect 134708 192976 134760 192982
rect 134708 192918 134760 192924
rect 134352 190426 134472 190454
rect 134248 148572 134300 148578
rect 134248 148514 134300 148520
rect 134444 148510 134472 190426
rect 135364 189854 135392 197474
rect 135456 194274 135484 199679
rect 135628 199650 135680 199656
rect 135536 199572 135588 199578
rect 135536 199514 135588 199520
rect 135548 199073 135576 199514
rect 135534 199064 135590 199073
rect 135534 198999 135590 199008
rect 135444 194268 135496 194274
rect 135444 194210 135496 194216
rect 135640 191162 135668 199650
rect 135732 191185 135760 199718
rect 135548 191134 135668 191162
rect 135718 191176 135774 191185
rect 135548 190126 135576 191134
rect 135718 191111 135774 191120
rect 135628 191072 135680 191078
rect 135628 191014 135680 191020
rect 135536 190120 135588 190126
rect 135536 190062 135588 190068
rect 135352 189848 135404 189854
rect 135352 189790 135404 189796
rect 134432 148504 134484 148510
rect 134432 148446 134484 148452
rect 135640 148170 135668 191014
rect 135824 189922 135852 199736
rect 135962 199730 135990 200124
rect 136054 199918 136082 200124
rect 136042 199912 136094 199918
rect 136042 199854 136094 199860
rect 136146 199730 136174 200124
rect 136238 199918 136266 200124
rect 136330 199918 136358 200124
rect 136226 199912 136278 199918
rect 136226 199854 136278 199860
rect 136318 199912 136370 199918
rect 136318 199854 136370 199860
rect 135962 199702 136036 199730
rect 135904 199640 135956 199646
rect 135904 199582 135956 199588
rect 135916 194206 135944 199582
rect 135904 194200 135956 194206
rect 135904 194142 135956 194148
rect 136008 191049 136036 199702
rect 136100 199702 136174 199730
rect 136272 199776 136324 199782
rect 136422 199764 136450 200124
rect 136514 199889 136542 200124
rect 136500 199880 136556 199889
rect 136500 199815 136556 199824
rect 136606 199764 136634 200124
rect 136272 199718 136324 199724
rect 136376 199736 136450 199764
rect 136560 199753 136634 199764
rect 136546 199744 136634 199753
rect 136100 194342 136128 199702
rect 136284 198734 136312 199718
rect 136192 198706 136312 198734
rect 136088 194336 136140 194342
rect 136088 194278 136140 194284
rect 136192 191078 136220 198706
rect 136376 194002 136404 199736
rect 136602 199736 136634 199744
rect 136698 199764 136726 200124
rect 136790 199889 136818 200124
rect 136882 199918 136910 200124
rect 136974 199918 137002 200124
rect 136870 199912 136922 199918
rect 136776 199880 136832 199889
rect 136870 199854 136922 199860
rect 136962 199912 137014 199918
rect 137066 199889 137094 200124
rect 137158 199918 137186 200124
rect 137146 199912 137198 199918
rect 136962 199854 137014 199860
rect 137052 199880 137108 199889
rect 136776 199815 136832 199824
rect 137146 199854 137198 199860
rect 137250 199850 137278 200124
rect 137052 199815 137108 199824
rect 137238 199844 137290 199850
rect 137238 199786 137290 199792
rect 136916 199776 136968 199782
rect 136698 199736 136772 199764
rect 136546 199679 136602 199688
rect 136640 199640 136692 199646
rect 136454 199608 136510 199617
rect 136638 199608 136640 199617
rect 136692 199608 136694 199617
rect 136454 199543 136510 199552
rect 136548 199572 136600 199578
rect 136468 199442 136496 199543
rect 136638 199543 136694 199552
rect 136548 199514 136600 199520
rect 136456 199436 136508 199442
rect 136456 199378 136508 199384
rect 136454 199064 136510 199073
rect 136454 198999 136510 199008
rect 136468 198354 136496 198999
rect 136560 198801 136588 199514
rect 136546 198792 136602 198801
rect 136546 198727 136602 198736
rect 136456 198348 136508 198354
rect 136456 198290 136508 198296
rect 136548 198348 136600 198354
rect 136548 198290 136600 198296
rect 136560 198121 136588 198290
rect 136546 198112 136602 198121
rect 136546 198047 136602 198056
rect 136640 197532 136692 197538
rect 136640 197474 136692 197480
rect 136364 193996 136416 194002
rect 136364 193938 136416 193944
rect 136652 193934 136680 197474
rect 136744 194546 136772 199736
rect 136822 199744 136878 199753
rect 136916 199718 136968 199724
rect 136822 199679 136878 199688
rect 136732 194540 136784 194546
rect 136732 194482 136784 194488
rect 136640 193928 136692 193934
rect 136640 193870 136692 193876
rect 136180 191072 136232 191078
rect 135994 191040 136050 191049
rect 136180 191014 136232 191020
rect 135994 190975 136050 190984
rect 136836 190454 136864 199679
rect 136928 194478 136956 199718
rect 137100 199708 137152 199714
rect 137100 199650 137152 199656
rect 137192 199708 137244 199714
rect 137342 199696 137370 200124
rect 137434 199918 137462 200124
rect 137526 199918 137554 200124
rect 137618 199918 137646 200124
rect 137422 199912 137474 199918
rect 137422 199854 137474 199860
rect 137514 199912 137566 199918
rect 137514 199854 137566 199860
rect 137606 199912 137658 199918
rect 137710 199889 137738 200124
rect 137606 199854 137658 199860
rect 137696 199880 137752 199889
rect 137696 199815 137752 199824
rect 137468 199776 137520 199782
rect 137468 199718 137520 199724
rect 137802 199730 137830 200124
rect 137894 199889 137922 200124
rect 137880 199880 137936 199889
rect 137880 199815 137936 199824
rect 137986 199730 138014 200124
rect 138078 199889 138106 200124
rect 138064 199880 138120 199889
rect 138064 199815 138120 199824
rect 138170 199730 138198 200124
rect 138262 199889 138290 200124
rect 138354 199918 138382 200124
rect 138342 199912 138394 199918
rect 138248 199880 138304 199889
rect 138446 199889 138474 200124
rect 138342 199854 138394 199860
rect 138432 199880 138488 199889
rect 138248 199815 138304 199824
rect 138432 199815 138488 199824
rect 138538 199764 138566 200124
rect 138630 199918 138658 200124
rect 138722 199918 138750 200124
rect 138814 199918 138842 200124
rect 138906 199918 138934 200124
rect 138618 199912 138670 199918
rect 138618 199854 138670 199860
rect 138710 199912 138762 199918
rect 138710 199854 138762 199860
rect 138802 199912 138854 199918
rect 138802 199854 138854 199860
rect 138894 199912 138946 199918
rect 138998 199889 139026 200124
rect 138894 199854 138946 199860
rect 138984 199880 139040 199889
rect 139090 199850 139118 200124
rect 138984 199815 139040 199824
rect 139078 199844 139130 199850
rect 139078 199786 139130 199792
rect 138848 199776 138900 199782
rect 138538 199736 138612 199764
rect 137342 199668 137416 199696
rect 137192 199650 137244 199656
rect 137112 195129 137140 199650
rect 137204 197538 137232 199650
rect 137284 199572 137336 199578
rect 137284 199514 137336 199520
rect 137192 197532 137244 197538
rect 137192 197474 137244 197480
rect 137296 195974 137324 199514
rect 137388 197985 137416 199668
rect 137374 197976 137430 197985
rect 137374 197911 137430 197920
rect 137296 195946 137416 195974
rect 137098 195120 137154 195129
rect 137098 195055 137154 195064
rect 136916 194472 136968 194478
rect 136916 194414 136968 194420
rect 136836 190426 137140 190454
rect 135812 189916 135864 189922
rect 135812 189858 135864 189864
rect 135628 148164 135680 148170
rect 135628 148106 135680 148112
rect 137112 147014 137140 190426
rect 137388 180794 137416 195946
rect 137480 193798 137508 199718
rect 137802 199702 137876 199730
rect 137986 199702 138060 199730
rect 138170 199702 138244 199730
rect 137652 199640 137704 199646
rect 137652 199582 137704 199588
rect 137560 199504 137612 199510
rect 137560 199446 137612 199452
rect 137572 198558 137600 199446
rect 137560 198552 137612 198558
rect 137560 198494 137612 198500
rect 137664 197849 137692 199582
rect 137744 198552 137796 198558
rect 137744 198494 137796 198500
rect 137650 197840 137706 197849
rect 137650 197775 137706 197784
rect 137756 196314 137784 198494
rect 137744 196308 137796 196314
rect 137744 196250 137796 196256
rect 137848 195974 137876 199702
rect 137928 199572 137980 199578
rect 137928 199514 137980 199520
rect 137664 195946 137876 195974
rect 137468 193792 137520 193798
rect 137468 193734 137520 193740
rect 137664 191214 137692 195946
rect 137652 191208 137704 191214
rect 137652 191150 137704 191156
rect 137940 183530 137968 199514
rect 138032 198558 138060 199702
rect 138110 199608 138166 199617
rect 138110 199543 138166 199552
rect 138020 198552 138072 198558
rect 138020 198494 138072 198500
rect 138020 198212 138072 198218
rect 138020 198154 138072 198160
rect 138032 194070 138060 198154
rect 138020 194064 138072 194070
rect 138020 194006 138072 194012
rect 138124 191350 138152 199543
rect 138112 191344 138164 191350
rect 138112 191286 138164 191292
rect 138216 190454 138244 199702
rect 138388 199640 138440 199646
rect 138294 199608 138350 199617
rect 138388 199582 138440 199588
rect 138294 199543 138350 199552
rect 138308 197198 138336 199543
rect 138296 197192 138348 197198
rect 138296 197134 138348 197140
rect 138400 191282 138428 199582
rect 138584 196897 138612 199736
rect 138848 199718 138900 199724
rect 138938 199744 138994 199753
rect 138664 199708 138716 199714
rect 138664 199650 138716 199656
rect 138756 199708 138808 199714
rect 138756 199650 138808 199656
rect 138570 196888 138626 196897
rect 138570 196823 138626 196832
rect 138388 191276 138440 191282
rect 138388 191218 138440 191224
rect 138676 191146 138704 199650
rect 138664 191140 138716 191146
rect 138664 191082 138716 191088
rect 138216 190426 138428 190454
rect 137928 183524 137980 183530
rect 137928 183466 137980 183472
rect 137296 180766 137416 180794
rect 137296 149705 137324 180766
rect 137282 149696 137338 149705
rect 137282 149631 137338 149640
rect 138400 148782 138428 190426
rect 138768 183297 138796 199650
rect 138860 197354 138888 199718
rect 139182 199730 139210 200124
rect 138938 199679 138994 199688
rect 139136 199702 139210 199730
rect 138952 198422 138980 199679
rect 139032 199572 139084 199578
rect 139032 199514 139084 199520
rect 139044 198966 139072 199514
rect 139032 198960 139084 198966
rect 139032 198902 139084 198908
rect 138940 198416 138992 198422
rect 138940 198358 138992 198364
rect 138860 197326 138980 197354
rect 138952 191418 138980 197326
rect 139136 191486 139164 199702
rect 139274 199696 139302 200124
rect 139366 199764 139394 200124
rect 139458 199923 139486 200124
rect 139444 199914 139500 199923
rect 139444 199849 139500 199858
rect 139366 199736 139440 199764
rect 139412 199730 139440 199736
rect 139412 199702 139486 199730
rect 139274 199668 139348 199696
rect 139320 199628 139348 199668
rect 139458 199628 139486 199702
rect 139550 199696 139578 200124
rect 139642 199764 139670 200124
rect 139734 199918 139762 200124
rect 139826 199918 139854 200124
rect 139918 199918 139946 200124
rect 140010 199918 140038 200124
rect 139722 199912 139774 199918
rect 139722 199854 139774 199860
rect 139814 199912 139866 199918
rect 139814 199854 139866 199860
rect 139906 199912 139958 199918
rect 139906 199854 139958 199860
rect 139998 199912 140050 199918
rect 140102 199889 140130 200124
rect 139998 199854 140050 199860
rect 140088 199880 140144 199889
rect 140088 199815 140144 199824
rect 140044 199776 140096 199782
rect 139642 199736 139716 199764
rect 139550 199668 139624 199696
rect 139320 199600 139394 199628
rect 139458 199617 139532 199628
rect 139458 199608 139546 199617
rect 139458 199600 139490 199608
rect 139216 199572 139268 199578
rect 139216 199514 139268 199520
rect 139228 197334 139256 199514
rect 139366 199458 139394 199600
rect 139490 199543 139546 199552
rect 139366 199430 139532 199458
rect 139400 199368 139452 199374
rect 139400 199310 139452 199316
rect 139306 199064 139362 199073
rect 139306 198999 139362 199008
rect 139216 197328 139268 197334
rect 139216 197270 139268 197276
rect 139320 195430 139348 198999
rect 139412 198121 139440 199310
rect 139504 198801 139532 199430
rect 139490 198792 139546 198801
rect 139490 198727 139546 198736
rect 139398 198112 139454 198121
rect 139398 198047 139454 198056
rect 139492 198008 139544 198014
rect 139492 197950 139544 197956
rect 139308 195424 139360 195430
rect 139308 195366 139360 195372
rect 139504 193186 139532 197950
rect 139492 193180 139544 193186
rect 139492 193122 139544 193128
rect 139124 191480 139176 191486
rect 139124 191422 139176 191428
rect 138940 191412 138992 191418
rect 138940 191354 138992 191360
rect 139596 190454 139624 199668
rect 139688 196790 139716 199736
rect 140044 199718 140096 199724
rect 139768 199708 139820 199714
rect 139768 199650 139820 199656
rect 139780 199374 139808 199650
rect 139952 199640 140004 199646
rect 139952 199582 140004 199588
rect 139964 199424 139992 199582
rect 139872 199396 139992 199424
rect 139768 199368 139820 199374
rect 139768 199310 139820 199316
rect 139872 198218 139900 199396
rect 139952 198960 140004 198966
rect 139952 198902 140004 198908
rect 139964 198665 139992 198902
rect 139950 198656 140006 198665
rect 139950 198591 140006 198600
rect 139860 198212 139912 198218
rect 139860 198154 139912 198160
rect 139858 198112 139914 198121
rect 139858 198047 139914 198056
rect 139676 196784 139728 196790
rect 139676 196726 139728 196732
rect 139872 192370 139900 198047
rect 139860 192364 139912 192370
rect 139860 192306 139912 192312
rect 140056 192302 140084 199718
rect 140194 199696 140222 200124
rect 140286 199918 140314 200124
rect 140274 199912 140326 199918
rect 140274 199854 140326 199860
rect 140148 199668 140222 199696
rect 140272 199710 140328 199719
rect 140148 198734 140176 199668
rect 140378 199696 140406 200124
rect 140470 199918 140498 200124
rect 140458 199912 140510 199918
rect 140458 199854 140510 199860
rect 140562 199730 140590 200124
rect 140654 199764 140682 200124
rect 140746 199918 140774 200124
rect 140734 199912 140786 199918
rect 140734 199854 140786 199860
rect 140654 199736 140728 199764
rect 140838 199753 140866 200124
rect 140516 199702 140590 199730
rect 140378 199668 140452 199696
rect 140272 199645 140328 199654
rect 140424 198734 140452 199668
rect 140148 198706 140268 198734
rect 140240 193866 140268 198706
rect 140332 198706 140452 198734
rect 140332 198121 140360 198706
rect 140318 198112 140374 198121
rect 140318 198047 140374 198056
rect 140516 198014 140544 199702
rect 140596 199640 140648 199646
rect 140596 199582 140648 199588
rect 140504 198008 140556 198014
rect 140504 197950 140556 197956
rect 140608 195974 140636 199582
rect 140700 199073 140728 199736
rect 140824 199744 140880 199753
rect 140824 199679 140880 199688
rect 140780 199640 140832 199646
rect 140780 199582 140832 199588
rect 140792 199510 140820 199582
rect 140930 199560 140958 200124
rect 141022 199889 141050 200124
rect 141008 199880 141064 199889
rect 141008 199815 141064 199824
rect 141114 199696 141142 200124
rect 141206 199918 141234 200124
rect 141194 199912 141246 199918
rect 141298 199889 141326 200124
rect 141194 199854 141246 199860
rect 141284 199880 141340 199889
rect 141284 199815 141340 199824
rect 141390 199764 141418 200124
rect 141482 199918 141510 200124
rect 141470 199912 141522 199918
rect 141574 199889 141602 200124
rect 141470 199854 141522 199860
rect 141560 199880 141616 199889
rect 141666 199850 141694 200124
rect 141560 199815 141616 199824
rect 141654 199844 141706 199850
rect 141654 199786 141706 199792
rect 141344 199736 141418 199764
rect 141514 199744 141570 199753
rect 141344 199730 141372 199736
rect 140884 199532 140958 199560
rect 141068 199668 141142 199696
rect 141252 199702 141372 199730
rect 140780 199504 140832 199510
rect 140780 199446 140832 199452
rect 140686 199064 140742 199073
rect 140686 198999 140742 199008
rect 140780 198076 140832 198082
rect 140780 198018 140832 198024
rect 140792 195974 140820 198018
rect 140884 197554 140912 199532
rect 140884 197526 141004 197554
rect 140516 195946 140636 195974
rect 140700 195946 140820 195974
rect 140516 195770 140544 195946
rect 140700 195838 140728 195946
rect 140688 195832 140740 195838
rect 140688 195774 140740 195780
rect 140504 195764 140556 195770
rect 140504 195706 140556 195712
rect 140228 193860 140280 193866
rect 140228 193802 140280 193808
rect 140044 192296 140096 192302
rect 140044 192238 140096 192244
rect 139596 190426 139808 190454
rect 138754 183288 138810 183297
rect 138754 183223 138810 183232
rect 138388 148776 138440 148782
rect 138388 148718 138440 148724
rect 139780 148442 139808 190426
rect 139768 148436 139820 148442
rect 139768 148378 139820 148384
rect 140976 148238 141004 197526
rect 141068 195702 141096 199668
rect 141148 199504 141200 199510
rect 141148 199446 141200 199452
rect 141160 198082 141188 199446
rect 141148 198076 141200 198082
rect 141148 198018 141200 198024
rect 141056 195696 141108 195702
rect 141056 195638 141108 195644
rect 141252 189990 141280 199702
rect 141758 199730 141786 200124
rect 141850 199918 141878 200124
rect 141942 199918 141970 200124
rect 141838 199912 141890 199918
rect 141838 199854 141890 199860
rect 141930 199912 141982 199918
rect 141930 199854 141982 199860
rect 141514 199679 141570 199688
rect 141608 199708 141660 199714
rect 141424 199640 141476 199646
rect 141330 199608 141386 199617
rect 141424 199582 141476 199588
rect 141330 199543 141386 199552
rect 141344 192681 141372 199543
rect 141330 192672 141386 192681
rect 141330 192607 141386 192616
rect 141240 189984 141292 189990
rect 141240 189926 141292 189932
rect 140964 148232 141016 148238
rect 140964 148174 141016 148180
rect 137100 147008 137152 147014
rect 137100 146950 137152 146956
rect 137008 144628 137060 144634
rect 137008 144570 137060 144576
rect 133144 143404 133196 143410
rect 133144 143346 133196 143352
rect 133156 139890 133184 143346
rect 135444 143336 135496 143342
rect 135444 143278 135496 143284
rect 134800 143268 134852 143274
rect 134800 143210 134852 143216
rect 134248 142928 134300 142934
rect 134248 142870 134300 142876
rect 133880 142248 133932 142254
rect 133880 142190 133932 142196
rect 133892 139890 133920 142190
rect 134260 139890 134288 142870
rect 134812 139890 134840 143210
rect 135456 139890 135484 143278
rect 136640 143200 136692 143206
rect 136640 143142 136692 143148
rect 135904 142792 135956 142798
rect 135904 142734 135956 142740
rect 135916 139890 135944 142734
rect 136652 139890 136680 143142
rect 137020 139890 137048 144570
rect 140870 144528 140926 144537
rect 140870 144463 140926 144472
rect 138662 143984 138718 143993
rect 138662 143919 138718 143928
rect 137560 143472 137612 143478
rect 137560 143414 137612 143420
rect 137572 139890 137600 143414
rect 138112 141704 138164 141710
rect 138112 141646 138164 141652
rect 138124 139890 138152 141646
rect 138676 139890 138704 143919
rect 139398 143848 139454 143857
rect 139398 143783 139454 143792
rect 139412 139890 139440 143783
rect 139768 143064 139820 143070
rect 139768 143006 139820 143012
rect 139780 139890 139808 143006
rect 140318 141808 140374 141817
rect 140318 141743 140374 141752
rect 140332 139890 140360 141743
rect 140884 139890 140912 144463
rect 141436 141137 141464 199582
rect 141528 198608 141556 199679
rect 141608 199650 141660 199656
rect 141712 199702 141786 199730
rect 141884 199776 141936 199782
rect 142034 199764 142062 200124
rect 142126 199923 142154 200124
rect 142112 199914 142168 199923
rect 142218 199918 142246 200124
rect 142112 199849 142168 199858
rect 142206 199912 142258 199918
rect 142206 199854 142258 199860
rect 141884 199718 141936 199724
rect 141988 199736 142062 199764
rect 142160 199776 142212 199782
rect 141620 198676 141648 199650
rect 141712 199628 141740 199702
rect 141712 199600 141832 199628
rect 141620 198648 141740 198676
rect 141528 198580 141648 198608
rect 141516 198484 141568 198490
rect 141516 198426 141568 198432
rect 141528 141273 141556 198426
rect 141620 192817 141648 198580
rect 141606 192808 141662 192817
rect 141606 192743 141662 192752
rect 141712 190194 141740 198648
rect 141700 190188 141752 190194
rect 141700 190130 141752 190136
rect 141804 188873 141832 199600
rect 141896 189786 141924 199718
rect 141988 196081 142016 199736
rect 142160 199718 142212 199724
rect 142068 199640 142120 199646
rect 142068 199582 142120 199588
rect 142080 198490 142108 199582
rect 142068 198484 142120 198490
rect 142068 198426 142120 198432
rect 142172 198336 142200 199718
rect 142310 199628 142338 200124
rect 142402 199918 142430 200124
rect 142494 199923 142522 200124
rect 142390 199912 142442 199918
rect 142390 199854 142442 199860
rect 142480 199914 142536 199923
rect 142480 199849 142536 199858
rect 142080 198308 142200 198336
rect 142264 199600 142338 199628
rect 142436 199640 142488 199646
rect 141974 196072 142030 196081
rect 141974 196007 142030 196016
rect 141974 195392 142030 195401
rect 141974 195327 142030 195336
rect 141988 195129 142016 195327
rect 141974 195120 142030 195129
rect 141974 195055 142030 195064
rect 142080 192642 142108 198308
rect 142264 196994 142292 199600
rect 142586 199628 142614 200124
rect 142678 199850 142706 200124
rect 142770 199918 142798 200124
rect 142758 199912 142810 199918
rect 142758 199854 142810 199860
rect 142666 199844 142718 199850
rect 142666 199786 142718 199792
rect 142862 199764 142890 200124
rect 142816 199736 142890 199764
rect 142712 199708 142764 199714
rect 142712 199650 142764 199656
rect 142586 199600 142660 199628
rect 142724 199617 142752 199650
rect 142436 199582 142488 199588
rect 142252 196988 142304 196994
rect 142252 196930 142304 196936
rect 142448 196042 142476 199582
rect 142436 196036 142488 196042
rect 142436 195978 142488 195984
rect 142632 192778 142660 199600
rect 142710 199608 142766 199617
rect 142710 199543 142766 199552
rect 142712 199504 142764 199510
rect 142712 199446 142764 199452
rect 142620 192772 142672 192778
rect 142620 192714 142672 192720
rect 142724 192658 142752 199446
rect 142068 192636 142120 192642
rect 142068 192578 142120 192584
rect 142540 192630 142752 192658
rect 141884 189780 141936 189786
rect 141884 189722 141936 189728
rect 141790 188864 141846 188873
rect 141790 188799 141846 188808
rect 142540 147082 142568 192630
rect 142816 192545 142844 199736
rect 142954 199696 142982 200124
rect 143046 199918 143074 200124
rect 143138 199918 143166 200124
rect 143034 199912 143086 199918
rect 143034 199854 143086 199860
rect 143126 199912 143178 199918
rect 143126 199854 143178 199860
rect 143230 199850 143258 200124
rect 143322 199918 143350 200124
rect 143310 199912 143362 199918
rect 143310 199854 143362 199860
rect 143218 199844 143270 199850
rect 143218 199786 143270 199792
rect 143170 199744 143226 199753
rect 142908 199668 142982 199696
rect 143080 199708 143132 199714
rect 142908 195974 142936 199668
rect 143414 199696 143442 200124
rect 143506 199889 143534 200124
rect 143492 199880 143548 199889
rect 143492 199815 143548 199824
rect 143598 199764 143626 200124
rect 143690 199918 143718 200124
rect 143678 199912 143730 199918
rect 143678 199854 143730 199860
rect 143170 199679 143226 199688
rect 143080 199650 143132 199656
rect 142988 199572 143040 199578
rect 142988 199514 143040 199520
rect 142896 195968 142948 195974
rect 142896 195910 142948 195916
rect 142802 192536 142858 192545
rect 142802 192471 142858 192480
rect 142620 191072 142672 191078
rect 142620 191014 142672 191020
rect 142632 149054 142660 191014
rect 143000 182174 143028 199514
rect 143092 195906 143120 199650
rect 143184 197266 143212 199679
rect 143368 199668 143442 199696
rect 143552 199736 143626 199764
rect 143264 199640 143316 199646
rect 143264 199582 143316 199588
rect 143172 197260 143224 197266
rect 143172 197202 143224 197208
rect 143080 195900 143132 195906
rect 143080 195842 143132 195848
rect 143276 191078 143304 199582
rect 143368 196518 143396 199668
rect 143448 199232 143500 199238
rect 143448 199174 143500 199180
rect 143460 199073 143488 199174
rect 143446 199064 143502 199073
rect 143446 198999 143502 199008
rect 143356 196512 143408 196518
rect 143356 196454 143408 196460
rect 143552 194177 143580 199736
rect 143782 199730 143810 200124
rect 143874 199918 143902 200124
rect 143966 199918 143994 200124
rect 143862 199912 143914 199918
rect 143862 199854 143914 199860
rect 143954 199912 144006 199918
rect 143954 199854 144006 199860
rect 143736 199702 143810 199730
rect 143908 199776 143960 199782
rect 144058 199764 144086 200124
rect 144150 199918 144178 200124
rect 144242 199918 144270 200124
rect 144138 199912 144190 199918
rect 144138 199854 144190 199860
rect 144230 199912 144282 199918
rect 144230 199854 144282 199860
rect 144334 199764 144362 200124
rect 143908 199718 143960 199724
rect 144012 199736 144086 199764
rect 144288 199736 144362 199764
rect 144426 199764 144454 200124
rect 144518 199923 144546 200124
rect 144504 199914 144560 199923
rect 144504 199849 144560 199858
rect 144610 199764 144638 200124
rect 144702 199918 144730 200124
rect 144690 199912 144742 199918
rect 144690 199854 144742 199860
rect 144426 199736 144500 199764
rect 144610 199736 144684 199764
rect 143632 199640 143684 199646
rect 143632 199582 143684 199588
rect 143644 198626 143672 199582
rect 143736 198762 143764 199702
rect 143816 199640 143868 199646
rect 143816 199582 143868 199588
rect 143724 198756 143776 198762
rect 143724 198698 143776 198704
rect 143632 198620 143684 198626
rect 143632 198562 143684 198568
rect 143828 197577 143856 199582
rect 143814 197568 143870 197577
rect 143814 197503 143870 197512
rect 143538 194168 143594 194177
rect 143538 194103 143594 194112
rect 143920 192846 143948 199718
rect 144012 197062 144040 199736
rect 144092 199640 144144 199646
rect 144092 199582 144144 199588
rect 144184 199640 144236 199646
rect 144184 199582 144236 199588
rect 144104 198937 144132 199582
rect 144196 198966 144224 199582
rect 144184 198960 144236 198966
rect 144090 198928 144146 198937
rect 144184 198902 144236 198908
rect 144090 198863 144146 198872
rect 144182 198792 144238 198801
rect 144092 198756 144144 198762
rect 144182 198727 144238 198736
rect 144092 198698 144144 198704
rect 144000 197056 144052 197062
rect 144000 196998 144052 197004
rect 144104 195634 144132 198698
rect 144092 195628 144144 195634
rect 144092 195570 144144 195576
rect 144090 195392 144146 195401
rect 144090 195327 144146 195336
rect 144104 195090 144132 195327
rect 144092 195084 144144 195090
rect 144092 195026 144144 195032
rect 143998 193216 144054 193225
rect 143998 193151 144054 193160
rect 144012 193118 144040 193151
rect 144000 193112 144052 193118
rect 144000 193054 144052 193060
rect 143908 192840 143960 192846
rect 143908 192782 143960 192788
rect 144196 192574 144224 198727
rect 144288 196858 144316 199736
rect 144472 198880 144500 199736
rect 144552 199640 144604 199646
rect 144552 199582 144604 199588
rect 144380 198852 144500 198880
rect 144380 198529 144408 198852
rect 144564 198830 144592 199582
rect 144552 198824 144604 198830
rect 144552 198766 144604 198772
rect 144366 198520 144422 198529
rect 144366 198455 144422 198464
rect 144552 197396 144604 197402
rect 144552 197338 144604 197344
rect 144276 196852 144328 196858
rect 144276 196794 144328 196800
rect 144184 192568 144236 192574
rect 144184 192510 144236 192516
rect 144564 192506 144592 197338
rect 144656 196382 144684 199736
rect 144794 199730 144822 200124
rect 144748 199702 144822 199730
rect 144644 196376 144696 196382
rect 144644 196318 144696 196324
rect 144748 195974 144776 199702
rect 144886 199628 144914 200124
rect 144978 199918 145006 200124
rect 144966 199912 145018 199918
rect 144966 199854 145018 199860
rect 145070 199628 145098 200124
rect 145162 199764 145190 200124
rect 145254 199918 145282 200124
rect 145242 199912 145294 199918
rect 145242 199854 145294 199860
rect 145346 199764 145374 200124
rect 145438 199923 145466 200124
rect 145424 199914 145480 199923
rect 145424 199849 145480 199858
rect 145530 199850 145558 200124
rect 145622 199850 145650 200124
rect 145714 199918 145742 200124
rect 145806 199918 145834 200124
rect 145898 199918 145926 200124
rect 145990 199918 146018 200124
rect 146082 199918 146110 200124
rect 145702 199912 145754 199918
rect 145702 199854 145754 199860
rect 145794 199912 145846 199918
rect 145794 199854 145846 199860
rect 145886 199912 145938 199918
rect 145886 199854 145938 199860
rect 145978 199912 146030 199918
rect 145978 199854 146030 199860
rect 146070 199912 146122 199918
rect 146174 199889 146202 200124
rect 146070 199854 146122 199860
rect 146160 199880 146216 199889
rect 145518 199844 145570 199850
rect 145518 199786 145570 199792
rect 145610 199844 145662 199850
rect 146160 199815 146216 199824
rect 145610 199786 145662 199792
rect 146116 199776 146168 199782
rect 145162 199736 145236 199764
rect 145346 199736 145420 199764
rect 144656 195946 144776 195974
rect 144840 199600 144914 199628
rect 145024 199600 145098 199628
rect 144552 192500 144604 192506
rect 144552 192442 144604 192448
rect 144656 192438 144684 195946
rect 144840 195158 144868 199600
rect 144920 199504 144972 199510
rect 144920 199446 144972 199452
rect 144932 197985 144960 199446
rect 144918 197976 144974 197985
rect 144918 197911 144974 197920
rect 145024 195566 145052 199600
rect 145104 199368 145156 199374
rect 145104 199310 145156 199316
rect 145116 197674 145144 199310
rect 145208 199306 145236 199736
rect 145288 199640 145340 199646
rect 145288 199582 145340 199588
rect 145196 199300 145248 199306
rect 145196 199242 145248 199248
rect 145300 197810 145328 199582
rect 145392 198393 145420 199736
rect 146266 199764 146294 200124
rect 146358 199918 146386 200124
rect 146346 199912 146398 199918
rect 146346 199854 146398 199860
rect 146450 199764 146478 200124
rect 146116 199718 146168 199724
rect 146220 199736 146294 199764
rect 146404 199736 146478 199764
rect 145472 199708 145524 199714
rect 145472 199650 145524 199656
rect 146024 199708 146076 199714
rect 146024 199650 146076 199656
rect 145378 198384 145434 198393
rect 145378 198319 145434 198328
rect 145288 197804 145340 197810
rect 145288 197746 145340 197752
rect 145104 197668 145156 197674
rect 145104 197610 145156 197616
rect 145484 196450 145512 199650
rect 145564 199640 145616 199646
rect 145564 199582 145616 199588
rect 145840 199640 145892 199646
rect 145840 199582 145892 199588
rect 145932 199640 145984 199646
rect 145932 199582 145984 199588
rect 145576 197849 145604 199582
rect 145656 199572 145708 199578
rect 145656 199514 145708 199520
rect 145668 199170 145696 199514
rect 145656 199164 145708 199170
rect 145656 199106 145708 199112
rect 145656 198552 145708 198558
rect 145656 198494 145708 198500
rect 145562 197840 145618 197849
rect 145562 197775 145618 197784
rect 145472 196444 145524 196450
rect 145472 196386 145524 196392
rect 145012 195560 145064 195566
rect 145012 195502 145064 195508
rect 144828 195152 144880 195158
rect 144828 195094 144880 195100
rect 145564 193248 145616 193254
rect 145564 193190 145616 193196
rect 144644 192432 144696 192438
rect 144644 192374 144696 192380
rect 143264 191072 143316 191078
rect 143264 191014 143316 191020
rect 143000 182146 143120 182174
rect 142620 149048 142672 149054
rect 142620 148990 142672 148996
rect 143092 148986 143120 182146
rect 143080 148980 143132 148986
rect 143080 148922 143132 148928
rect 142528 147076 142580 147082
rect 142528 147018 142580 147024
rect 144184 144560 144236 144566
rect 144184 144502 144236 144508
rect 142528 144492 142580 144498
rect 142528 144434 142580 144440
rect 141608 143132 141660 143138
rect 141608 143074 141660 143080
rect 141514 141264 141570 141273
rect 141514 141199 141570 141208
rect 141422 141128 141478 141137
rect 141422 141063 141478 141072
rect 141620 139890 141648 143074
rect 142250 141672 142306 141681
rect 142250 141607 142306 141616
rect 142264 139890 142292 141607
rect 142540 139890 142568 144434
rect 143080 142996 143132 143002
rect 143080 142938 143132 142944
rect 143092 139890 143120 142938
rect 143630 141536 143686 141545
rect 143630 141471 143686 141480
rect 143644 139890 143672 141471
rect 144196 139890 144224 144502
rect 145288 143608 145340 143614
rect 145288 143550 145340 143556
rect 145010 143168 145066 143177
rect 145010 143103 145066 143112
rect 145024 139890 145052 143103
rect 145300 139890 145328 143550
rect 145576 140350 145604 193190
rect 145668 148481 145696 198494
rect 145852 198354 145880 199582
rect 145840 198348 145892 198354
rect 145840 198290 145892 198296
rect 145944 197606 145972 199582
rect 146036 198150 146064 199650
rect 146024 198144 146076 198150
rect 146024 198086 146076 198092
rect 145932 197600 145984 197606
rect 145932 197542 145984 197548
rect 146128 195537 146156 199718
rect 146220 198694 146248 199736
rect 146404 199696 146432 199736
rect 146312 199668 146432 199696
rect 146542 199696 146570 200124
rect 146634 199764 146662 200124
rect 146726 199918 146754 200124
rect 146714 199912 146766 199918
rect 146714 199854 146766 199860
rect 146818 199764 146846 200124
rect 146634 199736 146708 199764
rect 146542 199668 146616 199696
rect 146208 198688 146260 198694
rect 146208 198630 146260 198636
rect 146114 195528 146170 195537
rect 146114 195463 146170 195472
rect 146312 194594 146340 199668
rect 146392 199572 146444 199578
rect 146392 199514 146444 199520
rect 146484 199572 146536 199578
rect 146484 199514 146536 199520
rect 146128 194566 146340 194594
rect 146128 193050 146156 194566
rect 146116 193044 146168 193050
rect 146116 192986 146168 192992
rect 145748 184748 145800 184754
rect 145748 184690 145800 184696
rect 145654 148472 145710 148481
rect 145654 148407 145710 148416
rect 145564 140344 145616 140350
rect 145564 140286 145616 140292
rect 133156 139862 133492 139890
rect 133892 139862 134044 139890
rect 134260 139862 134596 139890
rect 134812 139862 135148 139890
rect 135456 139862 135700 139890
rect 135916 139862 136252 139890
rect 136652 139862 136804 139890
rect 137020 139862 137356 139890
rect 137572 139862 137908 139890
rect 138124 139862 138460 139890
rect 138676 139862 139012 139890
rect 139412 139862 139564 139890
rect 139780 139862 140116 139890
rect 140332 139862 140668 139890
rect 140884 139862 141220 139890
rect 141620 139862 141772 139890
rect 142264 139862 142324 139890
rect 142540 139862 142876 139890
rect 143092 139862 143428 139890
rect 143644 139862 143980 139890
rect 144196 139862 144532 139890
rect 145024 139862 145084 139890
rect 145300 139862 145636 139890
rect 145760 139369 145788 184690
rect 146404 182174 146432 199514
rect 146496 197305 146524 199514
rect 146588 199034 146616 199668
rect 146576 199028 146628 199034
rect 146576 198970 146628 198976
rect 146680 197742 146708 199736
rect 146772 199736 146846 199764
rect 146772 197985 146800 199736
rect 146910 199696 146938 200124
rect 146864 199668 146938 199696
rect 146758 197976 146814 197985
rect 146758 197911 146814 197920
rect 146668 197736 146720 197742
rect 146668 197678 146720 197684
rect 146482 197296 146538 197305
rect 146482 197231 146538 197240
rect 146760 196036 146812 196042
rect 146760 195978 146812 195984
rect 146404 182146 146524 182174
rect 146496 146946 146524 182146
rect 146484 146940 146536 146946
rect 146484 146882 146536 146888
rect 146666 145888 146722 145897
rect 146666 145823 146722 145832
rect 146298 145752 146354 145761
rect 146298 145687 146354 145696
rect 145838 144392 145894 144401
rect 145838 144327 145894 144336
rect 145852 139890 145880 144327
rect 146312 143478 146340 145687
rect 146300 143472 146352 143478
rect 146300 143414 146352 143420
rect 146390 142896 146446 142905
rect 146390 142831 146446 142840
rect 146404 139890 146432 142831
rect 146680 140570 146708 145823
rect 146772 140690 146800 195978
rect 146864 195809 146892 199668
rect 147002 199628 147030 200124
rect 146956 199600 147030 199628
rect 146956 197402 146984 199600
rect 147094 199560 147122 200124
rect 147186 199918 147214 200124
rect 147278 199918 147306 200124
rect 147370 199918 147398 200124
rect 147174 199912 147226 199918
rect 147174 199854 147226 199860
rect 147266 199912 147318 199918
rect 147266 199854 147318 199860
rect 147358 199912 147410 199918
rect 147358 199854 147410 199860
rect 147220 199776 147272 199782
rect 147462 199764 147490 200124
rect 147554 199923 147582 200124
rect 147540 199914 147596 199923
rect 147540 199849 147596 199858
rect 147646 199764 147674 200124
rect 147738 199918 147766 200124
rect 147726 199912 147778 199918
rect 147830 199889 147858 200124
rect 147726 199854 147778 199860
rect 147816 199880 147872 199889
rect 147922 199850 147950 200124
rect 148014 199923 148042 200124
rect 148000 199914 148056 199923
rect 148106 199918 148134 200124
rect 148198 199923 148226 200124
rect 147816 199815 147872 199824
rect 147910 199844 147962 199850
rect 148000 199849 148056 199858
rect 148094 199912 148146 199918
rect 148094 199854 148146 199860
rect 148184 199914 148240 199923
rect 148290 199918 148318 200124
rect 148382 199918 148410 200124
rect 148184 199849 148240 199858
rect 148278 199912 148330 199918
rect 148278 199854 148330 199860
rect 148370 199912 148422 199918
rect 148370 199854 148422 199860
rect 147910 199786 147962 199792
rect 148474 199764 148502 200124
rect 148566 199918 148594 200124
rect 148554 199912 148606 199918
rect 148554 199854 148606 199860
rect 147220 199718 147272 199724
rect 147416 199736 147490 199764
rect 147600 199736 147674 199764
rect 148428 199753 148502 199764
rect 148554 199776 148606 199782
rect 148414 199744 148502 199753
rect 147048 199532 147122 199560
rect 147048 199073 147076 199532
rect 147034 199064 147090 199073
rect 147034 198999 147090 199008
rect 147232 198937 147260 199718
rect 147312 199708 147364 199714
rect 147312 199650 147364 199656
rect 147218 198928 147274 198937
rect 147218 198863 147274 198872
rect 147218 198792 147274 198801
rect 147218 198727 147274 198736
rect 146944 197396 146996 197402
rect 146944 197338 146996 197344
rect 147036 197396 147088 197402
rect 147036 197338 147088 197344
rect 146850 195800 146906 195809
rect 146850 195735 146906 195744
rect 147048 191834 147076 197338
rect 146864 191806 147076 191834
rect 146864 141642 146892 191806
rect 147232 180794 147260 198727
rect 147324 197402 147352 199650
rect 147312 197396 147364 197402
rect 147312 197338 147364 197344
rect 147416 196042 147444 199736
rect 147600 199102 147628 199736
rect 147772 199708 147824 199714
rect 147772 199650 147824 199656
rect 148048 199708 148100 199714
rect 148048 199650 148100 199656
rect 148232 199708 148284 199714
rect 148232 199650 148284 199656
rect 148324 199708 148376 199714
rect 148470 199736 148502 199744
rect 148552 199744 148554 199753
rect 148606 199744 148608 199753
rect 148414 199679 148470 199688
rect 148552 199679 148608 199688
rect 148324 199650 148376 199656
rect 147678 199608 147734 199617
rect 147678 199543 147734 199552
rect 147588 199096 147640 199102
rect 147588 199038 147640 199044
rect 147692 198422 147720 199543
rect 147680 198416 147732 198422
rect 147680 198358 147732 198364
rect 147404 196036 147456 196042
rect 147404 195978 147456 195984
rect 147784 190454 147812 199650
rect 147954 198928 148010 198937
rect 147954 198863 147956 198872
rect 148008 198863 148010 198872
rect 147956 198834 148008 198840
rect 148060 197946 148088 199650
rect 148140 199436 148192 199442
rect 148140 199378 148192 199384
rect 148152 198937 148180 199378
rect 148138 198928 148194 198937
rect 148138 198863 148194 198872
rect 148048 197940 148100 197946
rect 148048 197882 148100 197888
rect 148244 193662 148272 199650
rect 148336 195226 148364 199650
rect 148658 199628 148686 200124
rect 148750 199753 148778 200124
rect 148842 199764 148870 200124
rect 148934 199918 148962 200124
rect 148922 199912 148974 199918
rect 148922 199854 148974 199860
rect 149026 199764 149054 200124
rect 148736 199744 148792 199753
rect 148842 199736 148916 199764
rect 148736 199679 148792 199688
rect 148784 199640 148836 199646
rect 148414 199608 148470 199617
rect 148658 199600 148732 199628
rect 148414 199543 148470 199552
rect 148324 195220 148376 195226
rect 148324 195162 148376 195168
rect 148232 193656 148284 193662
rect 148232 193598 148284 193604
rect 147784 190426 147904 190454
rect 147588 189168 147640 189174
rect 147588 189110 147640 189116
rect 146956 180766 147260 180794
rect 146852 141636 146904 141642
rect 146852 141578 146904 141584
rect 146956 140758 146984 180766
rect 147600 147121 147628 189110
rect 147586 147112 147642 147121
rect 147586 147047 147642 147056
rect 147876 145654 147904 190426
rect 148048 184952 148100 184958
rect 148048 184894 148100 184900
rect 148060 151814 148088 184894
rect 148428 182174 148456 199543
rect 148508 198620 148560 198626
rect 148508 198562 148560 198568
rect 148520 198286 148548 198562
rect 148508 198280 148560 198286
rect 148508 198222 148560 198228
rect 148704 191834 148732 199600
rect 148782 199608 148784 199617
rect 148836 199608 148838 199617
rect 148782 199543 148838 199552
rect 148612 191806 148732 191834
rect 148612 191185 148640 191806
rect 148598 191176 148654 191185
rect 148598 191111 148654 191120
rect 148600 185836 148652 185842
rect 148600 185778 148652 185784
rect 147968 151786 148088 151814
rect 148244 182146 148456 182174
rect 147864 145648 147916 145654
rect 147678 145616 147734 145625
rect 147864 145590 147916 145596
rect 147678 145551 147734 145560
rect 146944 140752 146996 140758
rect 146944 140694 146996 140700
rect 146760 140684 146812 140690
rect 146760 140626 146812 140632
rect 146680 140542 146892 140570
rect 146864 139890 146892 140542
rect 147692 139890 147720 145551
rect 147968 140282 147996 151786
rect 148046 143032 148102 143041
rect 148046 142967 148102 142976
rect 147956 140276 148008 140282
rect 147956 140218 148008 140224
rect 148060 139890 148088 142967
rect 148244 140418 148272 182146
rect 148612 180794 148640 185778
rect 148888 184958 148916 199736
rect 148980 199736 149054 199764
rect 148980 199646 149008 199736
rect 149118 199696 149146 200124
rect 149210 199730 149238 200124
rect 149302 199918 149330 200124
rect 149394 199923 149422 200124
rect 149290 199912 149342 199918
rect 149290 199854 149342 199860
rect 149380 199914 149436 199923
rect 149486 199918 149514 200124
rect 149578 199918 149606 200124
rect 149670 199923 149698 200124
rect 149380 199849 149436 199858
rect 149474 199912 149526 199918
rect 149474 199854 149526 199860
rect 149566 199912 149618 199918
rect 149566 199854 149618 199860
rect 149656 199914 149712 199923
rect 149656 199849 149712 199858
rect 149762 199730 149790 200124
rect 149854 199918 149882 200124
rect 149842 199912 149894 199918
rect 149946 199889 149974 200124
rect 150038 199918 150066 200124
rect 150026 199912 150078 199918
rect 149842 199854 149894 199860
rect 149932 199880 149988 199889
rect 150026 199854 150078 199860
rect 149932 199815 149988 199824
rect 149210 199702 149468 199730
rect 149072 199668 149146 199696
rect 148968 199640 149020 199646
rect 148968 199582 149020 199588
rect 149072 199578 149100 199668
rect 149244 199640 149296 199646
rect 149244 199582 149296 199588
rect 149060 199572 149112 199578
rect 149060 199514 149112 199520
rect 149152 199572 149204 199578
rect 149152 199514 149204 199520
rect 148968 199504 149020 199510
rect 148966 199472 148968 199481
rect 149020 199472 149022 199481
rect 148966 199407 149022 199416
rect 149164 191834 149192 199514
rect 149072 191806 149192 191834
rect 148968 191548 149020 191554
rect 148968 191490 149020 191496
rect 148876 184952 148928 184958
rect 148876 184894 148928 184900
rect 148336 180766 148640 180794
rect 148336 148306 148364 180766
rect 148324 148300 148376 148306
rect 148324 148242 148376 148248
rect 148600 146940 148652 146946
rect 148600 146882 148652 146888
rect 148232 140412 148284 140418
rect 148232 140354 148284 140360
rect 148612 139890 148640 146882
rect 148980 145654 149008 191490
rect 149072 191049 149100 191806
rect 149058 191040 149114 191049
rect 149058 190975 149114 190984
rect 149256 149734 149284 199582
rect 149440 198626 149468 199702
rect 149520 199708 149572 199714
rect 149520 199650 149572 199656
rect 149716 199702 149790 199730
rect 149888 199776 149940 199782
rect 149888 199718 149940 199724
rect 149428 198620 149480 198626
rect 149428 198562 149480 198568
rect 149426 198520 149482 198529
rect 149426 198455 149482 198464
rect 149244 149728 149296 149734
rect 149244 149670 149296 149676
rect 148968 145648 149020 145654
rect 148968 145590 149020 145596
rect 149152 143472 149204 143478
rect 149152 143414 149204 143420
rect 149164 139890 149192 143414
rect 149440 140214 149468 198455
rect 149532 194041 149560 199650
rect 149610 199472 149666 199481
rect 149610 199407 149666 199416
rect 149518 194032 149574 194041
rect 149518 193967 149574 193976
rect 149624 193254 149652 199407
rect 149612 193248 149664 193254
rect 149612 193190 149664 193196
rect 149716 193032 149744 199702
rect 149796 199640 149848 199646
rect 149796 199582 149848 199588
rect 149808 196489 149836 199582
rect 149900 199209 149928 199718
rect 150130 199696 150158 200124
rect 149992 199668 150158 199696
rect 149886 199200 149942 199209
rect 149886 199135 149942 199144
rect 149992 196926 150020 199668
rect 150222 199628 150250 200124
rect 150314 199714 150342 200124
rect 150302 199708 150354 199714
rect 150406 199696 150434 200124
rect 150498 199918 150526 200124
rect 150590 199918 150618 200124
rect 150682 199918 150710 200124
rect 150774 199923 150802 200124
rect 150486 199912 150538 199918
rect 150486 199854 150538 199860
rect 150578 199912 150630 199918
rect 150578 199854 150630 199860
rect 150670 199912 150722 199918
rect 150670 199854 150722 199860
rect 150760 199914 150816 199923
rect 150866 199918 150894 200124
rect 150958 199918 150986 200124
rect 151050 199918 151078 200124
rect 150760 199849 150816 199858
rect 150854 199912 150906 199918
rect 150854 199854 150906 199860
rect 150946 199912 150998 199918
rect 150946 199854 150998 199860
rect 151038 199912 151090 199918
rect 151038 199854 151090 199860
rect 150900 199776 150952 199782
rect 151142 199764 151170 200124
rect 151234 199889 151262 200124
rect 151220 199880 151276 199889
rect 151220 199815 151276 199824
rect 151326 199764 151354 200124
rect 151418 199889 151446 200124
rect 151404 199880 151460 199889
rect 151404 199815 151460 199824
rect 151510 199764 151538 200124
rect 151142 199736 151216 199764
rect 151326 199736 151400 199764
rect 150900 199718 150952 199724
rect 150406 199668 150480 199696
rect 150302 199650 150354 199656
rect 150176 199600 150250 199628
rect 150072 199572 150124 199578
rect 150072 199514 150124 199520
rect 150084 197033 150112 199514
rect 150070 197024 150126 197033
rect 150070 196959 150126 196968
rect 149980 196920 150032 196926
rect 149980 196862 150032 196868
rect 149794 196480 149850 196489
rect 149794 196415 149850 196424
rect 149624 193004 149744 193032
rect 149624 192914 149652 193004
rect 149612 192908 149664 192914
rect 149612 192850 149664 192856
rect 149704 192228 149756 192234
rect 149704 192170 149756 192176
rect 149716 145790 149744 192170
rect 149796 183252 149848 183258
rect 149796 183194 149848 183200
rect 149808 148850 149836 183194
rect 150176 180794 150204 199600
rect 150348 199572 150400 199578
rect 150348 199514 150400 199520
rect 150360 195673 150388 199514
rect 150452 199345 150480 199668
rect 150808 199640 150860 199646
rect 150808 199582 150860 199588
rect 150532 199504 150584 199510
rect 150532 199446 150584 199452
rect 150438 199336 150494 199345
rect 150438 199271 150494 199280
rect 150346 195664 150402 195673
rect 150346 195599 150402 195608
rect 150544 192710 150572 199446
rect 150716 199436 150768 199442
rect 150716 199378 150768 199384
rect 150532 192704 150584 192710
rect 150532 192646 150584 192652
rect 150728 192506 150756 199378
rect 150820 195673 150848 199582
rect 150912 199458 150940 199718
rect 151084 199640 151136 199646
rect 151084 199582 151136 199588
rect 150912 199430 151032 199458
rect 150900 199368 150952 199374
rect 150900 199310 150952 199316
rect 150806 195664 150862 195673
rect 150806 195599 150862 195608
rect 150716 192500 150768 192506
rect 150716 192442 150768 192448
rect 150624 191276 150676 191282
rect 150624 191218 150676 191224
rect 150084 180766 150204 180794
rect 149796 148844 149848 148850
rect 149796 148786 149848 148792
rect 149704 145784 149756 145790
rect 149704 145726 149756 145732
rect 149702 142760 149758 142769
rect 149702 142695 149758 142704
rect 149428 140208 149480 140214
rect 149428 140150 149480 140156
rect 149716 139890 149744 142695
rect 150084 140146 150112 180766
rect 150636 146985 150664 191218
rect 150622 146976 150678 146985
rect 150622 146911 150678 146920
rect 150438 141400 150494 141409
rect 150438 141335 150494 141344
rect 150072 140140 150124 140146
rect 150072 140082 150124 140088
rect 150452 139890 150480 141335
rect 145852 139862 146188 139890
rect 146404 139862 146740 139890
rect 146864 139862 147292 139890
rect 147692 139862 147844 139890
rect 148060 139862 148396 139890
rect 148612 139862 148948 139890
rect 149164 139862 149500 139890
rect 149716 139862 150052 139890
rect 150452 139862 150604 139890
rect 150912 139369 150940 199310
rect 151004 199102 151032 199430
rect 150992 199096 151044 199102
rect 150992 199038 151044 199044
rect 151096 196586 151124 199582
rect 151188 199458 151216 199736
rect 151188 199430 151308 199458
rect 151176 199368 151228 199374
rect 151176 199310 151228 199316
rect 151084 196580 151136 196586
rect 151084 196522 151136 196528
rect 151188 183258 151216 199310
rect 151280 196081 151308 199430
rect 151266 196072 151322 196081
rect 151266 196007 151322 196016
rect 151372 191834 151400 199736
rect 151464 199736 151538 199764
rect 151602 199764 151630 200124
rect 151694 199918 151722 200124
rect 151682 199912 151734 199918
rect 151682 199854 151734 199860
rect 151786 199764 151814 200124
rect 151878 199918 151906 200124
rect 151970 199918 151998 200124
rect 151866 199912 151918 199918
rect 151866 199854 151918 199860
rect 151958 199912 152010 199918
rect 152062 199889 152090 200124
rect 151958 199854 152010 199860
rect 152048 199880 152104 199889
rect 152048 199815 152104 199824
rect 151602 199736 151676 199764
rect 151464 197878 151492 199736
rect 151544 199640 151596 199646
rect 151544 199582 151596 199588
rect 151556 199306 151584 199582
rect 151544 199300 151596 199306
rect 151544 199242 151596 199248
rect 151452 197872 151504 197878
rect 151452 197814 151504 197820
rect 151648 191834 151676 199736
rect 151740 199736 151814 199764
rect 151912 199776 151964 199782
rect 151740 199481 151768 199736
rect 152154 199764 152182 200124
rect 151912 199718 151964 199724
rect 152108 199736 152182 199764
rect 151726 199472 151782 199481
rect 151726 199407 151782 199416
rect 151728 198280 151780 198286
rect 151728 198222 151780 198228
rect 151280 191806 151400 191834
rect 151556 191806 151676 191834
rect 151280 190454 151308 191806
rect 151556 191282 151584 191806
rect 151544 191276 151596 191282
rect 151544 191218 151596 191224
rect 151280 190426 151492 190454
rect 151176 183252 151228 183258
rect 151176 183194 151228 183200
rect 151464 145858 151492 190426
rect 151740 149705 151768 198222
rect 151924 197354 151952 199718
rect 152004 199708 152056 199714
rect 152004 199650 152056 199656
rect 151832 197326 151952 197354
rect 151832 192234 151860 197326
rect 152016 197169 152044 199650
rect 152002 197160 152058 197169
rect 152002 197095 152058 197104
rect 151820 192228 151872 192234
rect 151820 192170 151872 192176
rect 152108 149802 152136 199736
rect 152246 199696 152274 200124
rect 152338 199918 152366 200124
rect 152430 199918 152458 200124
rect 152522 199923 152550 200124
rect 152326 199912 152378 199918
rect 152326 199854 152378 199860
rect 152418 199912 152470 199918
rect 152418 199854 152470 199860
rect 152508 199914 152564 199923
rect 152508 199849 152564 199858
rect 152200 199668 152274 199696
rect 152464 199708 152516 199714
rect 152200 183569 152228 199668
rect 152614 199696 152642 200124
rect 152706 199918 152734 200124
rect 152798 199923 152826 200124
rect 152694 199912 152746 199918
rect 152694 199854 152746 199860
rect 152784 199914 152840 199923
rect 152890 199918 152918 200124
rect 152784 199849 152840 199858
rect 152878 199912 152930 199918
rect 152878 199854 152930 199860
rect 152982 199850 153010 200124
rect 153074 199923 153102 200124
rect 153060 199914 153116 199923
rect 153166 199918 153194 200124
rect 153258 199918 153286 200124
rect 152970 199844 153022 199850
rect 153060 199849 153116 199858
rect 153154 199912 153206 199918
rect 153154 199854 153206 199860
rect 153246 199912 153298 199918
rect 153246 199854 153298 199860
rect 152970 199786 153022 199792
rect 152924 199708 152976 199714
rect 152614 199668 152688 199696
rect 152464 199650 152516 199656
rect 152476 187694 152504 199650
rect 152660 196625 152688 199668
rect 152924 199650 152976 199656
rect 153016 199708 153068 199714
rect 153350 199696 153378 200124
rect 153442 199918 153470 200124
rect 153430 199912 153482 199918
rect 153430 199854 153482 199860
rect 153534 199764 153562 200124
rect 153626 199889 153654 200124
rect 153718 199918 153746 200124
rect 153706 199912 153758 199918
rect 153612 199880 153668 199889
rect 153706 199854 153758 199860
rect 153612 199815 153668 199824
rect 153016 199650 153068 199656
rect 153304 199668 153378 199696
rect 153488 199736 153562 199764
rect 153660 199776 153712 199782
rect 152832 199572 152884 199578
rect 152832 199514 152884 199520
rect 152646 196616 152702 196625
rect 152646 196551 152702 196560
rect 152384 187666 152504 187694
rect 152844 187694 152872 199514
rect 152936 195362 152964 199650
rect 152924 195356 152976 195362
rect 152924 195298 152976 195304
rect 152844 187666 152964 187694
rect 152186 183560 152242 183569
rect 152186 183495 152242 183504
rect 152096 149796 152148 149802
rect 152096 149738 152148 149744
rect 151726 149696 151782 149705
rect 151726 149631 151782 149640
rect 151452 145852 151504 145858
rect 151452 145794 151504 145800
rect 151912 144356 151964 144362
rect 151912 144298 151964 144304
rect 150990 144120 151046 144129
rect 150990 144055 151046 144064
rect 151004 139890 151032 144055
rect 151360 142860 151412 142866
rect 151360 142802 151412 142808
rect 151372 139890 151400 142802
rect 151924 139890 151952 144298
rect 152384 141574 152412 187666
rect 152556 185700 152608 185706
rect 152556 185642 152608 185648
rect 152464 144424 152516 144430
rect 152464 144366 152516 144372
rect 152372 141568 152424 141574
rect 152372 141510 152424 141516
rect 152476 139890 152504 144366
rect 152568 144265 152596 185642
rect 152936 182174 152964 187666
rect 153028 185706 153056 199650
rect 153304 193050 153332 199668
rect 153384 199572 153436 199578
rect 153384 199514 153436 199520
rect 153396 197742 153424 199514
rect 153488 198734 153516 199736
rect 153810 199764 153838 200124
rect 153902 199918 153930 200124
rect 153890 199912 153942 199918
rect 153890 199854 153942 199860
rect 153994 199764 154022 200124
rect 154086 199850 154114 200124
rect 154178 199889 154206 200124
rect 154270 199918 154298 200124
rect 154362 199918 154390 200124
rect 154258 199912 154310 199918
rect 154164 199880 154220 199889
rect 154074 199844 154126 199850
rect 154258 199854 154310 199860
rect 154350 199912 154402 199918
rect 154454 199889 154482 200124
rect 154350 199854 154402 199860
rect 154440 199880 154496 199889
rect 154164 199815 154220 199824
rect 154440 199815 154496 199824
rect 154074 199786 154126 199792
rect 153660 199718 153712 199724
rect 153764 199736 153838 199764
rect 153948 199736 154022 199764
rect 154212 199776 154264 199782
rect 153672 199034 153700 199718
rect 153660 199028 153712 199034
rect 153660 198970 153712 198976
rect 153488 198706 153608 198734
rect 153384 197736 153436 197742
rect 153384 197678 153436 197684
rect 153292 193044 153344 193050
rect 153292 192986 153344 192992
rect 153292 191208 153344 191214
rect 153292 191150 153344 191156
rect 153016 185700 153068 185706
rect 153016 185642 153068 185648
rect 152936 182146 153056 182174
rect 153028 145722 153056 182146
rect 153016 145716 153068 145722
rect 153016 145658 153068 145664
rect 152554 144256 152610 144265
rect 152554 144191 152610 144200
rect 153304 141506 153332 191150
rect 153384 185496 153436 185502
rect 153384 185438 153436 185444
rect 153396 148918 153424 185438
rect 153580 182174 153608 198706
rect 153658 197432 153714 197441
rect 153658 197367 153714 197376
rect 153672 190913 153700 197367
rect 153658 190904 153714 190913
rect 153658 190839 153714 190848
rect 153488 182146 153608 182174
rect 153764 182174 153792 199736
rect 153844 199640 153896 199646
rect 153844 199582 153896 199588
rect 153856 189417 153884 199582
rect 153948 198966 153976 199736
rect 154546 199764 154574 200124
rect 154212 199718 154264 199724
rect 154500 199736 154574 199764
rect 154028 199640 154080 199646
rect 154080 199600 154160 199628
rect 154028 199582 154080 199588
rect 154026 199336 154082 199345
rect 154026 199271 154082 199280
rect 153936 198960 153988 198966
rect 153936 198902 153988 198908
rect 154040 191321 154068 199271
rect 154026 191312 154082 191321
rect 154026 191247 154082 191256
rect 153842 189408 153898 189417
rect 153842 189343 153898 189352
rect 154132 185502 154160 199600
rect 154224 195634 154252 199718
rect 154304 199640 154356 199646
rect 154304 199582 154356 199588
rect 154212 195628 154264 195634
rect 154212 195570 154264 195576
rect 154316 191214 154344 199582
rect 154500 199442 154528 199736
rect 154638 199696 154666 200124
rect 154730 199764 154758 200124
rect 154822 199889 154850 200124
rect 154808 199880 154864 199889
rect 154808 199815 154864 199824
rect 154914 199764 154942 200124
rect 154730 199736 154804 199764
rect 154592 199668 154666 199696
rect 154488 199436 154540 199442
rect 154488 199378 154540 199384
rect 154396 199300 154448 199306
rect 154396 199242 154448 199248
rect 154408 193118 154436 199242
rect 154592 198734 154620 199668
rect 154672 199572 154724 199578
rect 154672 199514 154724 199520
rect 154684 199186 154712 199514
rect 154776 199306 154804 199736
rect 154868 199736 154942 199764
rect 154868 199646 154896 199736
rect 155006 199730 155034 200124
rect 155098 199918 155126 200124
rect 155086 199912 155138 199918
rect 155086 199854 155138 199860
rect 155190 199764 155218 200124
rect 155282 199923 155310 200124
rect 155268 199914 155324 199923
rect 155374 199918 155402 200124
rect 155268 199849 155324 199858
rect 155362 199912 155414 199918
rect 155362 199854 155414 199860
rect 155144 199736 155218 199764
rect 155316 199776 155368 199782
rect 155006 199702 155080 199730
rect 154856 199640 154908 199646
rect 154856 199582 154908 199588
rect 154856 199504 154908 199510
rect 154854 199472 154856 199481
rect 154908 199472 154910 199481
rect 154854 199407 154910 199416
rect 154856 199368 154908 199374
rect 154856 199310 154908 199316
rect 154946 199336 155002 199345
rect 154764 199300 154816 199306
rect 154764 199242 154816 199248
rect 154684 199158 154804 199186
rect 154592 198706 154712 198734
rect 154578 198656 154634 198665
rect 154578 198591 154634 198600
rect 154592 198393 154620 198591
rect 154578 198384 154634 198393
rect 154578 198319 154634 198328
rect 154396 193112 154448 193118
rect 154396 193054 154448 193060
rect 154304 191208 154356 191214
rect 154304 191150 154356 191156
rect 154684 185842 154712 198706
rect 154776 189174 154804 199158
rect 154868 195401 154896 199310
rect 154946 199271 155002 199280
rect 154960 198665 154988 199271
rect 154946 198656 155002 198665
rect 154946 198591 155002 198600
rect 154854 195392 154910 195401
rect 154854 195327 154910 195336
rect 155052 194041 155080 199702
rect 155038 194032 155094 194041
rect 155038 193967 155094 193976
rect 154764 189168 154816 189174
rect 154764 189110 154816 189116
rect 155144 187694 155172 199736
rect 155316 199718 155368 199724
rect 155466 199730 155494 200124
rect 155558 199918 155586 200124
rect 155650 199918 155678 200124
rect 155546 199912 155598 199918
rect 155546 199854 155598 199860
rect 155638 199912 155690 199918
rect 155638 199854 155690 199860
rect 155592 199776 155644 199782
rect 155328 199238 155356 199718
rect 155466 199702 155540 199730
rect 155742 199764 155770 200124
rect 155834 199889 155862 200124
rect 155820 199880 155876 199889
rect 155820 199815 155876 199824
rect 155592 199718 155644 199724
rect 155696 199736 155770 199764
rect 155926 199764 155954 200124
rect 156018 199918 156046 200124
rect 156110 199918 156138 200124
rect 156202 199918 156230 200124
rect 156006 199912 156058 199918
rect 156006 199854 156058 199860
rect 156098 199912 156150 199918
rect 156098 199854 156150 199860
rect 156190 199912 156242 199918
rect 156190 199854 156242 199860
rect 156294 199850 156322 200124
rect 156386 199918 156414 200124
rect 156374 199912 156426 199918
rect 156374 199854 156426 199860
rect 156282 199844 156334 199850
rect 156282 199786 156334 199792
rect 156144 199776 156196 199782
rect 155926 199736 156000 199764
rect 155408 199572 155460 199578
rect 155408 199514 155460 199520
rect 155316 199232 155368 199238
rect 155316 199174 155368 199180
rect 155420 197946 155448 199514
rect 155408 197940 155460 197946
rect 155408 197882 155460 197888
rect 155052 187666 155172 187694
rect 154856 187604 154908 187610
rect 154856 187546 154908 187552
rect 154672 185836 154724 185842
rect 154672 185778 154724 185784
rect 154764 185632 154816 185638
rect 154764 185574 154816 185580
rect 154120 185496 154172 185502
rect 154120 185438 154172 185444
rect 153764 182146 154068 182174
rect 153384 148912 153436 148918
rect 153384 148854 153436 148860
rect 153488 148714 153516 182146
rect 153476 148708 153528 148714
rect 153476 148650 153528 148656
rect 153658 142216 153714 142225
rect 153658 142151 153714 142160
rect 153292 141500 153344 141506
rect 153292 141442 153344 141448
rect 153672 139890 153700 142151
rect 153752 141432 153804 141438
rect 153752 141374 153804 141380
rect 151004 139862 151156 139890
rect 151372 139862 151708 139890
rect 151924 139862 152260 139890
rect 152476 139862 152812 139890
rect 153364 139862 153700 139890
rect 153764 139890 153792 141374
rect 153764 139862 153916 139890
rect 154040 139369 154068 182146
rect 154488 144356 154540 144362
rect 154488 144298 154540 144304
rect 154500 140162 154528 144298
rect 154454 140134 154528 140162
rect 154454 139876 154482 140134
rect 154776 140049 154804 185574
rect 154868 149841 154896 187546
rect 155052 182174 155080 187666
rect 155512 185638 155540 199702
rect 155500 185632 155552 185638
rect 155500 185574 155552 185580
rect 155604 182174 155632 199718
rect 155696 187610 155724 199736
rect 155868 199640 155920 199646
rect 155868 199582 155920 199588
rect 155774 199336 155830 199345
rect 155774 199271 155830 199280
rect 155684 187604 155736 187610
rect 155684 187546 155736 187552
rect 155052 182146 155172 182174
rect 155604 182146 155724 182174
rect 155144 180794 155172 182146
rect 155052 180766 155172 180794
rect 155052 150113 155080 180766
rect 155038 150104 155094 150113
rect 155038 150039 155094 150048
rect 154854 149832 154910 149841
rect 154854 149767 154910 149776
rect 155314 142760 155370 142769
rect 155314 142695 155370 142704
rect 154762 140040 154818 140049
rect 154762 139975 154818 139984
rect 155328 139890 155356 142695
rect 155592 142248 155644 142254
rect 155592 142190 155644 142196
rect 155604 140162 155632 142190
rect 155020 139862 155356 139890
rect 155558 140134 155632 140162
rect 155558 139876 155586 140134
rect 155696 139369 155724 182146
rect 155788 151814 155816 199271
rect 155880 199170 155908 199582
rect 155868 199164 155920 199170
rect 155868 199106 155920 199112
rect 155972 198082 156000 199736
rect 156478 199764 156506 200124
rect 156144 199718 156196 199724
rect 156432 199736 156506 199764
rect 156052 199708 156104 199714
rect 156052 199650 156104 199656
rect 155960 198076 156012 198082
rect 155960 198018 156012 198024
rect 156064 195906 156092 199650
rect 156052 195900 156104 195906
rect 156052 195842 156104 195848
rect 156156 194954 156184 199718
rect 156236 199708 156288 199714
rect 156236 199650 156288 199656
rect 156328 199708 156380 199714
rect 156328 199650 156380 199656
rect 156144 194948 156196 194954
rect 156144 194890 156196 194896
rect 156248 184754 156276 199650
rect 156340 192574 156368 199650
rect 156432 198354 156460 199736
rect 156570 199696 156598 200124
rect 156662 199918 156690 200124
rect 156650 199912 156702 199918
rect 156650 199854 156702 199860
rect 156754 199764 156782 200124
rect 156524 199668 156598 199696
rect 156708 199736 156782 199764
rect 156420 198348 156472 198354
rect 156420 198290 156472 198296
rect 156524 198121 156552 199668
rect 156708 199424 156736 199736
rect 156846 199696 156874 200124
rect 156938 199764 156966 200124
rect 157030 199923 157058 200124
rect 157016 199914 157072 199923
rect 157016 199849 157072 199858
rect 156938 199736 157012 199764
rect 156616 199396 156736 199424
rect 156800 199668 156874 199696
rect 156510 198112 156566 198121
rect 156510 198047 156566 198056
rect 156616 195430 156644 199396
rect 156800 198734 156828 199668
rect 156984 199481 157012 199736
rect 157122 199696 157150 200124
rect 157076 199668 157150 199696
rect 156970 199472 157026 199481
rect 156880 199436 156932 199442
rect 156970 199407 157026 199416
rect 156880 199378 156932 199384
rect 156892 198937 156920 199378
rect 156972 199300 157024 199306
rect 156972 199242 157024 199248
rect 156878 198928 156934 198937
rect 156878 198863 156934 198872
rect 156984 198801 157012 199242
rect 156708 198706 156828 198734
rect 156970 198792 157026 198801
rect 156970 198727 157026 198736
rect 156708 198558 156736 198706
rect 156788 198620 156840 198626
rect 156788 198562 156840 198568
rect 156696 198552 156748 198558
rect 156696 198494 156748 198500
rect 156604 195424 156656 195430
rect 156604 195366 156656 195372
rect 156800 195022 156828 198562
rect 157076 198506 157104 199668
rect 157214 199628 157242 200124
rect 157168 199600 157242 199628
rect 157168 199442 157196 199600
rect 157306 199560 157334 200124
rect 157398 199918 157426 200124
rect 157386 199912 157438 199918
rect 157386 199854 157438 199860
rect 157386 199776 157438 199782
rect 157386 199718 157438 199724
rect 157490 199730 157518 200124
rect 157582 199918 157610 200124
rect 157570 199912 157622 199918
rect 157570 199854 157622 199860
rect 157674 199764 157702 200124
rect 157766 199918 157794 200124
rect 157858 199918 157886 200124
rect 157950 199918 157978 200124
rect 158042 199918 158070 200124
rect 157754 199912 157806 199918
rect 157754 199854 157806 199860
rect 157846 199912 157898 199918
rect 157846 199854 157898 199860
rect 157938 199912 157990 199918
rect 157938 199854 157990 199860
rect 158030 199912 158082 199918
rect 158030 199854 158082 199860
rect 158134 199764 158162 200124
rect 158226 199918 158254 200124
rect 158318 199918 158346 200124
rect 158214 199912 158266 199918
rect 158214 199854 158266 199860
rect 158306 199912 158358 199918
rect 158306 199854 158358 199860
rect 158410 199764 158438 200124
rect 158502 199918 158530 200124
rect 158490 199912 158542 199918
rect 158490 199854 158542 199860
rect 157628 199736 157702 199764
rect 158088 199736 158162 199764
rect 158272 199736 158438 199764
rect 157398 199628 157426 199718
rect 157490 199702 157564 199730
rect 157398 199600 157472 199628
rect 157306 199532 157380 199560
rect 157156 199436 157208 199442
rect 157156 199378 157208 199384
rect 157248 199368 157300 199374
rect 157154 199336 157210 199345
rect 157248 199310 157300 199316
rect 157154 199271 157210 199280
rect 157168 198626 157196 199271
rect 157260 198830 157288 199310
rect 157248 198824 157300 198830
rect 157248 198766 157300 198772
rect 157156 198620 157208 198626
rect 157156 198562 157208 198568
rect 156984 198478 157104 198506
rect 156788 195016 156840 195022
rect 156788 194958 156840 194964
rect 156328 192568 156380 192574
rect 156328 192510 156380 192516
rect 156236 184748 156288 184754
rect 156236 184690 156288 184696
rect 156984 180794 157012 198478
rect 157064 198416 157116 198422
rect 157064 198358 157116 198364
rect 156524 180766 157012 180794
rect 155788 151786 155908 151814
rect 155880 139369 155908 151786
rect 156418 144256 156474 144265
rect 156418 144191 156474 144200
rect 156432 139890 156460 144191
rect 156524 140185 156552 180766
rect 156970 142896 157026 142905
rect 156970 142831 157026 142840
rect 156510 140176 156566 140185
rect 156510 140111 156566 140120
rect 156984 139890 157012 142831
rect 156124 139862 156460 139890
rect 156676 139862 157012 139890
rect 157076 139369 157104 198358
rect 157156 195900 157208 195906
rect 157156 195842 157208 195848
rect 157168 149977 157196 195842
rect 157352 195265 157380 199532
rect 157444 198422 157472 199600
rect 157432 198416 157484 198422
rect 157432 198358 157484 198364
rect 157430 198248 157486 198257
rect 157430 198183 157486 198192
rect 157444 197713 157472 198183
rect 157430 197704 157486 197713
rect 157430 197639 157486 197648
rect 157536 196897 157564 199702
rect 157522 196888 157578 196897
rect 157522 196823 157578 196832
rect 157338 195256 157394 195265
rect 157338 195191 157394 195200
rect 157628 191554 157656 199736
rect 157800 199708 157852 199714
rect 157800 199650 157852 199656
rect 157708 199640 157760 199646
rect 157708 199582 157760 199588
rect 157720 196761 157748 199582
rect 157812 198490 157840 199650
rect 157892 199572 157944 199578
rect 157892 199514 157944 199520
rect 157904 198801 157932 199514
rect 157984 199504 158036 199510
rect 157984 199446 158036 199452
rect 157890 198792 157946 198801
rect 157890 198727 157946 198736
rect 157800 198484 157852 198490
rect 157800 198426 157852 198432
rect 157996 197354 158024 199446
rect 158088 198422 158116 199736
rect 158168 199640 158220 199646
rect 158168 199582 158220 199588
rect 158076 198416 158128 198422
rect 158076 198358 158128 198364
rect 157904 197326 158024 197354
rect 157706 196752 157762 196761
rect 157706 196687 157762 196696
rect 157616 191548 157668 191554
rect 157616 191490 157668 191496
rect 157904 180794 157932 197326
rect 158180 195974 158208 199582
rect 158272 199209 158300 199736
rect 158444 199640 158496 199646
rect 158594 199628 158622 200124
rect 158686 199918 158714 200124
rect 158778 199918 158806 200124
rect 158870 199918 158898 200124
rect 158674 199912 158726 199918
rect 158674 199854 158726 199860
rect 158766 199912 158818 199918
rect 158766 199854 158818 199860
rect 158858 199912 158910 199918
rect 158858 199854 158910 199860
rect 158720 199776 158772 199782
rect 158720 199718 158772 199724
rect 158812 199776 158864 199782
rect 158812 199718 158864 199724
rect 158444 199582 158496 199588
rect 158548 199600 158622 199628
rect 158352 199572 158404 199578
rect 158352 199514 158404 199520
rect 158258 199200 158314 199209
rect 158258 199135 158314 199144
rect 158364 198734 158392 199514
rect 158272 198706 158392 198734
rect 158272 198257 158300 198706
rect 158258 198248 158314 198257
rect 158258 198183 158314 198192
rect 158180 195946 158300 195974
rect 158076 195288 158128 195294
rect 158076 195230 158128 195236
rect 157444 180766 157932 180794
rect 157154 149968 157210 149977
rect 157154 149903 157210 149912
rect 157444 147393 157472 180766
rect 157430 147384 157486 147393
rect 157430 147319 157486 147328
rect 158088 145761 158116 195230
rect 158272 190454 158300 195946
rect 158456 195294 158484 199582
rect 158548 199345 158576 199600
rect 158628 199504 158680 199510
rect 158628 199446 158680 199452
rect 158534 199336 158590 199345
rect 158534 199271 158590 199280
rect 158534 199200 158590 199209
rect 158534 199135 158590 199144
rect 158548 199102 158576 199135
rect 158536 199096 158588 199102
rect 158536 199038 158588 199044
rect 158640 195566 158668 199446
rect 158732 198286 158760 199718
rect 158720 198280 158772 198286
rect 158720 198222 158772 198228
rect 158824 195673 158852 199718
rect 158962 199696 158990 200124
rect 159054 199764 159082 200124
rect 159146 199918 159174 200124
rect 159134 199912 159186 199918
rect 159134 199854 159186 199860
rect 159054 199736 159128 199764
rect 158962 199668 159036 199696
rect 158904 199572 158956 199578
rect 158904 199514 158956 199520
rect 158916 199481 158944 199514
rect 158902 199472 158958 199481
rect 158902 199407 158958 199416
rect 159008 199034 159036 199668
rect 158996 199028 159048 199034
rect 158996 198970 159048 198976
rect 159100 198734 159128 199736
rect 159238 199696 159266 200124
rect 159330 199918 159358 200124
rect 159318 199912 159370 199918
rect 159318 199854 159370 199860
rect 159422 199764 159450 200124
rect 159514 199918 159542 200124
rect 159502 199912 159554 199918
rect 159502 199854 159554 199860
rect 159606 199782 159634 200124
rect 159698 199850 159726 200124
rect 159790 199850 159818 200124
rect 159882 199850 159910 200124
rect 159974 199918 160002 200124
rect 160066 199918 160094 200124
rect 160158 199918 160186 200124
rect 159962 199912 160014 199918
rect 159962 199854 160014 199860
rect 160054 199912 160106 199918
rect 160054 199854 160106 199860
rect 160146 199912 160198 199918
rect 160250 199889 160278 200124
rect 160146 199854 160198 199860
rect 160236 199880 160292 199889
rect 159686 199844 159738 199850
rect 159686 199786 159738 199792
rect 159778 199844 159830 199850
rect 159778 199786 159830 199792
rect 159870 199844 159922 199850
rect 160236 199815 160292 199824
rect 159870 199786 159922 199792
rect 159594 199776 159646 199782
rect 159422 199736 159496 199764
rect 159238 199668 159312 199696
rect 159180 199572 159232 199578
rect 159180 199514 159232 199520
rect 159008 198706 159128 198734
rect 158904 195968 158956 195974
rect 158904 195910 158956 195916
rect 158810 195664 158866 195673
rect 158810 195599 158866 195608
rect 158628 195560 158680 195566
rect 158628 195502 158680 195508
rect 158812 195356 158864 195362
rect 158812 195298 158864 195304
rect 158444 195288 158496 195294
rect 158444 195230 158496 195236
rect 158272 190426 158576 190454
rect 158548 150249 158576 190426
rect 158534 150240 158590 150249
rect 158824 150210 158852 195298
rect 158916 150278 158944 195910
rect 159008 150346 159036 198706
rect 159192 197577 159220 199514
rect 159284 199442 159312 199668
rect 159364 199640 159416 199646
rect 159364 199582 159416 199588
rect 159272 199436 159324 199442
rect 159272 199378 159324 199384
rect 159178 197568 159234 197577
rect 159178 197503 159234 197512
rect 159088 195696 159140 195702
rect 159088 195638 159140 195644
rect 158996 150340 159048 150346
rect 158996 150282 159048 150288
rect 158904 150272 158956 150278
rect 158904 150214 158956 150220
rect 158534 150175 158590 150184
rect 158812 150204 158864 150210
rect 158812 150146 158864 150152
rect 159100 149666 159128 195638
rect 159376 195362 159404 199582
rect 159468 196625 159496 199736
rect 159962 199776 160014 199782
rect 159594 199718 159646 199724
rect 159928 199724 159962 199730
rect 159928 199718 160014 199724
rect 160192 199776 160244 199782
rect 160192 199718 160244 199724
rect 159732 199708 159784 199714
rect 159732 199650 159784 199656
rect 159824 199708 159876 199714
rect 159824 199650 159876 199656
rect 159928 199702 160002 199718
rect 159548 199640 159600 199646
rect 159548 199582 159600 199588
rect 159454 196616 159510 196625
rect 159454 196551 159510 196560
rect 159560 195702 159588 199582
rect 159640 199436 159692 199442
rect 159640 199378 159692 199384
rect 159652 197810 159680 199378
rect 159640 197804 159692 197810
rect 159640 197746 159692 197752
rect 159744 196761 159772 199650
rect 159730 196752 159786 196761
rect 159730 196687 159786 196696
rect 159836 195974 159864 199650
rect 159824 195968 159876 195974
rect 159824 195910 159876 195916
rect 159548 195696 159600 195702
rect 159548 195638 159600 195644
rect 159364 195356 159416 195362
rect 159364 195298 159416 195304
rect 159928 193214 159956 199702
rect 160008 199572 160060 199578
rect 160008 199514 160060 199520
rect 160100 199572 160152 199578
rect 160100 199514 160152 199520
rect 160020 199238 160048 199514
rect 160008 199232 160060 199238
rect 160008 199174 160060 199180
rect 160112 197418 160140 199514
rect 160204 198734 160232 199718
rect 160342 199696 160370 200124
rect 160434 199764 160462 200124
rect 160526 199918 160554 200124
rect 160514 199912 160566 199918
rect 160514 199854 160566 199860
rect 160618 199850 160646 200124
rect 160606 199844 160658 199850
rect 160606 199786 160658 199792
rect 160434 199736 160508 199764
rect 160342 199668 160416 199696
rect 160204 198706 160324 198734
rect 160112 197390 160232 197418
rect 160100 197328 160152 197334
rect 160100 197270 160152 197276
rect 160008 196444 160060 196450
rect 160008 196386 160060 196392
rect 159560 193186 159956 193214
rect 159088 149660 159140 149666
rect 159088 149602 159140 149608
rect 158074 145752 158130 145761
rect 158074 145687 158130 145696
rect 159456 144424 159508 144430
rect 159456 144366 159508 144372
rect 158074 144120 158130 144129
rect 158074 144055 158130 144064
rect 157340 142248 157392 142254
rect 157340 142190 157392 142196
rect 157352 142118 157380 142190
rect 157340 142112 157392 142118
rect 157340 142054 157392 142060
rect 157156 141432 157208 141438
rect 157156 141374 157208 141380
rect 157168 139890 157196 141374
rect 158088 139890 158116 144055
rect 158628 142860 158680 142866
rect 158628 142802 158680 142808
rect 158640 139890 158668 142802
rect 159180 142248 159232 142254
rect 159180 142190 159232 142196
rect 159192 139890 159220 142190
rect 159468 140162 159496 144366
rect 157168 139862 157228 139890
rect 157780 139862 158116 139890
rect 158332 139862 158668 139890
rect 158884 139862 159220 139890
rect 159422 140134 159496 140162
rect 159422 139876 159450 140134
rect 159560 139369 159588 193186
rect 160020 180794 160048 196386
rect 159744 180766 160048 180794
rect 159744 139369 159772 180766
rect 160112 144566 160140 197270
rect 160204 195537 160232 197390
rect 160190 195528 160246 195537
rect 160190 195463 160246 195472
rect 160192 185428 160244 185434
rect 160192 185370 160244 185376
rect 160204 145790 160232 185370
rect 160296 150414 160324 198706
rect 160388 196314 160416 199668
rect 160376 196308 160428 196314
rect 160376 196250 160428 196256
rect 160376 196104 160428 196110
rect 160376 196046 160428 196052
rect 160388 152998 160416 196046
rect 160480 153134 160508 199736
rect 160710 199628 160738 200124
rect 160802 199918 160830 200124
rect 160894 199918 160922 200124
rect 160986 199918 161014 200124
rect 161078 199918 161106 200124
rect 160790 199912 160842 199918
rect 160790 199854 160842 199860
rect 160882 199912 160934 199918
rect 160882 199854 160934 199860
rect 160974 199912 161026 199918
rect 160974 199854 161026 199860
rect 161066 199912 161118 199918
rect 161066 199854 161118 199860
rect 160836 199776 160888 199782
rect 160836 199718 160888 199724
rect 160928 199776 160980 199782
rect 161170 199764 161198 200124
rect 160928 199718 160980 199724
rect 161124 199736 161198 199764
rect 160664 199600 160738 199628
rect 160560 199504 160612 199510
rect 160560 199446 160612 199452
rect 160572 186930 160600 199446
rect 160560 186924 160612 186930
rect 160560 186866 160612 186872
rect 160664 185434 160692 199600
rect 160744 199504 160796 199510
rect 160744 199446 160796 199452
rect 160756 190505 160784 199446
rect 160848 196178 160876 199718
rect 160836 196172 160888 196178
rect 160836 196114 160888 196120
rect 160940 196110 160968 199718
rect 161020 199708 161072 199714
rect 161020 199650 161072 199656
rect 161032 197305 161060 199650
rect 161018 197296 161074 197305
rect 161018 197231 161074 197240
rect 161124 196246 161152 199736
rect 161262 199696 161290 200124
rect 161354 199918 161382 200124
rect 161446 199918 161474 200124
rect 161342 199912 161394 199918
rect 161342 199854 161394 199860
rect 161434 199912 161486 199918
rect 161434 199854 161486 199860
rect 161538 199850 161566 200124
rect 161526 199844 161578 199850
rect 161526 199786 161578 199792
rect 161216 199668 161290 199696
rect 161388 199708 161440 199714
rect 161216 197334 161244 199668
rect 161388 199650 161440 199656
rect 161296 199572 161348 199578
rect 161296 199514 161348 199520
rect 161308 197441 161336 199514
rect 161294 197432 161350 197441
rect 161294 197367 161350 197376
rect 161204 197328 161256 197334
rect 161204 197270 161256 197276
rect 161400 196858 161428 199650
rect 161480 199640 161532 199646
rect 161480 199582 161532 199588
rect 161492 197538 161520 199582
rect 161630 199560 161658 200124
rect 161722 199918 161750 200124
rect 161710 199912 161762 199918
rect 161710 199854 161762 199860
rect 161814 199764 161842 200124
rect 161906 199889 161934 200124
rect 161998 199918 162026 200124
rect 161986 199912 162038 199918
rect 161892 199880 161948 199889
rect 161986 199854 162038 199860
rect 161892 199815 161948 199824
rect 162090 199764 162118 200124
rect 161768 199736 161842 199764
rect 162044 199736 162118 199764
rect 161630 199532 161704 199560
rect 161572 199436 161624 199442
rect 161572 199378 161624 199384
rect 161480 197532 161532 197538
rect 161480 197474 161532 197480
rect 161480 197396 161532 197402
rect 161480 197338 161532 197344
rect 161388 196852 161440 196858
rect 161388 196794 161440 196800
rect 161112 196240 161164 196246
rect 161112 196182 161164 196188
rect 160928 196104 160980 196110
rect 160928 196046 160980 196052
rect 160742 190496 160798 190505
rect 160742 190431 160798 190440
rect 161386 190360 161442 190369
rect 161386 190295 161442 190304
rect 160652 185428 160704 185434
rect 160652 185370 160704 185376
rect 161400 180849 161428 190295
rect 161386 180840 161442 180849
rect 161386 180775 161442 180784
rect 161386 180704 161442 180713
rect 161386 180639 161442 180648
rect 161400 171193 161428 180639
rect 161386 171184 161442 171193
rect 161386 171119 161442 171128
rect 161386 171048 161442 171057
rect 161386 170983 161442 170992
rect 161400 161537 161428 170983
rect 161386 161528 161442 161537
rect 161386 161463 161442 161472
rect 161386 161392 161442 161401
rect 161386 161327 161442 161336
rect 160468 153128 160520 153134
rect 160468 153070 160520 153076
rect 160376 152992 160428 152998
rect 160376 152934 160428 152940
rect 161400 151881 161428 161327
rect 161386 151872 161442 151881
rect 161386 151807 161442 151816
rect 161386 151736 161442 151745
rect 161386 151671 161442 151680
rect 160284 150408 160336 150414
rect 160284 150350 160336 150356
rect 160192 145784 160244 145790
rect 160192 145726 160244 145732
rect 160652 145716 160704 145722
rect 160652 145658 160704 145664
rect 160100 144560 160152 144566
rect 160100 144502 160152 144508
rect 160558 144392 160614 144401
rect 160558 144327 160614 144336
rect 160006 143032 160062 143041
rect 160006 142967 160062 142976
rect 160020 140162 160048 142967
rect 160572 140162 160600 144327
rect 159974 140134 160048 140162
rect 160526 140134 160600 140162
rect 159974 139876 160002 140134
rect 160526 139876 160554 140134
rect 160664 139890 160692 145658
rect 161400 142361 161428 151671
rect 161492 148986 161520 197338
rect 161584 153066 161612 199378
rect 161676 198393 161704 199532
rect 161768 199442 161796 199736
rect 161940 199708 161992 199714
rect 161940 199650 161992 199656
rect 161848 199572 161900 199578
rect 161848 199514 161900 199520
rect 161756 199436 161808 199442
rect 161756 199378 161808 199384
rect 161662 198384 161718 198393
rect 161662 198319 161718 198328
rect 161756 197532 161808 197538
rect 161756 197474 161808 197480
rect 161664 196716 161716 196722
rect 161664 196658 161716 196664
rect 161572 153060 161624 153066
rect 161572 153002 161624 153008
rect 161676 152425 161704 196658
rect 161768 153202 161796 197474
rect 161860 196654 161888 199514
rect 161952 196994 161980 199650
rect 162044 197402 162072 199736
rect 162182 199696 162210 200124
rect 162136 199668 162210 199696
rect 162136 199345 162164 199668
rect 162274 199628 162302 200124
rect 162366 199918 162394 200124
rect 162458 199918 162486 200124
rect 162550 199918 162578 200124
rect 162354 199912 162406 199918
rect 162354 199854 162406 199860
rect 162446 199912 162498 199918
rect 162446 199854 162498 199860
rect 162538 199912 162590 199918
rect 162642 199889 162670 200124
rect 162734 199918 162762 200124
rect 162826 199918 162854 200124
rect 162918 199918 162946 200124
rect 162722 199912 162774 199918
rect 162538 199854 162590 199860
rect 162628 199880 162684 199889
rect 162722 199854 162774 199860
rect 162814 199912 162866 199918
rect 162814 199854 162866 199860
rect 162906 199912 162958 199918
rect 162906 199854 162958 199860
rect 162628 199815 162684 199824
rect 162676 199776 162728 199782
rect 162228 199600 162302 199628
rect 162504 199724 162676 199730
rect 162504 199718 162728 199724
rect 162768 199776 162820 199782
rect 162768 199718 162820 199724
rect 162860 199776 162912 199782
rect 163010 199764 163038 200124
rect 162860 199718 162912 199724
rect 162964 199736 163038 199764
rect 163102 199764 163130 200124
rect 163194 199918 163222 200124
rect 163286 199918 163314 200124
rect 163182 199912 163234 199918
rect 163182 199854 163234 199860
rect 163274 199912 163326 199918
rect 163274 199854 163326 199860
rect 163378 199764 163406 200124
rect 163470 199889 163498 200124
rect 163562 199918 163590 200124
rect 163654 199918 163682 200124
rect 163746 199918 163774 200124
rect 163550 199912 163602 199918
rect 163456 199880 163512 199889
rect 163550 199854 163602 199860
rect 163642 199912 163694 199918
rect 163642 199854 163694 199860
rect 163734 199912 163786 199918
rect 163838 199889 163866 200124
rect 163734 199854 163786 199860
rect 163824 199880 163880 199889
rect 163456 199815 163512 199824
rect 163824 199815 163880 199824
rect 163102 199736 163176 199764
rect 163378 199736 163452 199764
rect 162504 199702 162716 199718
rect 162122 199336 162178 199345
rect 162122 199271 162178 199280
rect 162032 197396 162084 197402
rect 162032 197338 162084 197344
rect 162228 197198 162256 199600
rect 162400 199572 162452 199578
rect 162400 199514 162452 199520
rect 162308 199504 162360 199510
rect 162308 199446 162360 199452
rect 162320 199102 162348 199446
rect 162308 199096 162360 199102
rect 162308 199038 162360 199044
rect 162216 197192 162268 197198
rect 162216 197134 162268 197140
rect 161940 196988 161992 196994
rect 161940 196930 161992 196936
rect 162412 196722 162440 199514
rect 162504 196761 162532 199702
rect 162584 199640 162636 199646
rect 162584 199582 162636 199588
rect 162490 196752 162546 196761
rect 162400 196716 162452 196722
rect 162490 196687 162546 196696
rect 162400 196658 162452 196664
rect 161848 196648 161900 196654
rect 161848 196590 161900 196596
rect 162596 195430 162624 199582
rect 162676 199436 162728 199442
rect 162676 199378 162728 199384
rect 162688 197470 162716 199378
rect 162676 197464 162728 197470
rect 162676 197406 162728 197412
rect 162780 196160 162808 199718
rect 162872 199442 162900 199718
rect 162860 199436 162912 199442
rect 162860 199378 162912 199384
rect 162964 197402 162992 199736
rect 163044 199504 163096 199510
rect 163044 199446 163096 199452
rect 163056 197577 163084 199446
rect 163148 199102 163176 199736
rect 163228 199708 163280 199714
rect 163228 199650 163280 199656
rect 163136 199096 163188 199102
rect 163136 199038 163188 199044
rect 163042 197568 163098 197577
rect 163042 197503 163098 197512
rect 163044 197464 163096 197470
rect 163044 197406 163096 197412
rect 162952 197396 163004 197402
rect 162952 197338 163004 197344
rect 162860 197056 162912 197062
rect 162860 196998 162912 197004
rect 162688 196132 162808 196160
rect 162688 195770 162716 196132
rect 162768 196036 162820 196042
rect 162768 195978 162820 195984
rect 162676 195764 162728 195770
rect 162676 195706 162728 195712
rect 162584 195424 162636 195430
rect 162584 195366 162636 195372
rect 161756 153196 161808 153202
rect 161756 153138 161808 153144
rect 162780 152522 162808 195978
rect 162768 152516 162820 152522
rect 162768 152458 162820 152464
rect 161662 152416 161718 152425
rect 161662 152351 161718 152360
rect 161480 148980 161532 148986
rect 161480 148922 161532 148928
rect 162766 144528 162822 144537
rect 162492 144492 162544 144498
rect 162766 144463 162822 144472
rect 162492 144434 162544 144440
rect 161938 143304 161994 143313
rect 161938 143239 161994 143248
rect 161386 142352 161442 142361
rect 161386 142287 161442 142296
rect 161480 142248 161532 142254
rect 161480 142190 161532 142196
rect 161492 142089 161520 142190
rect 161478 142080 161534 142089
rect 161478 142015 161534 142024
rect 161952 139890 161980 143239
rect 162504 139890 162532 144434
rect 162780 140162 162808 144463
rect 162872 141409 162900 196998
rect 162950 191176 163006 191185
rect 162950 191111 163006 191120
rect 162964 148646 162992 191111
rect 163056 152930 163084 197406
rect 163136 182436 163188 182442
rect 163136 182378 163188 182384
rect 163044 152924 163096 152930
rect 163044 152866 163096 152872
rect 163148 152561 163176 182378
rect 163134 152552 163190 152561
rect 163134 152487 163190 152496
rect 163240 152454 163268 199650
rect 163320 199640 163372 199646
rect 163320 199582 163372 199588
rect 163424 199594 163452 199736
rect 163930 199730 163958 200124
rect 164022 199918 164050 200124
rect 164010 199912 164062 199918
rect 164010 199854 164062 199860
rect 164114 199764 164142 200124
rect 164206 199918 164234 200124
rect 164194 199912 164246 199918
rect 164194 199854 164246 199860
rect 164114 199736 164188 199764
rect 163596 199708 163648 199714
rect 163930 199702 164004 199730
rect 163596 199650 163648 199656
rect 163332 199424 163360 199582
rect 163424 199566 163544 199594
rect 163332 199396 163452 199424
rect 163424 197441 163452 199396
rect 163410 197432 163466 197441
rect 163320 197396 163372 197402
rect 163410 197367 163466 197376
rect 163320 197338 163372 197344
rect 163332 193186 163360 197338
rect 163516 197130 163544 199566
rect 163504 197124 163556 197130
rect 163504 197066 163556 197072
rect 163320 193180 163372 193186
rect 163320 193122 163372 193128
rect 163608 189417 163636 199650
rect 163688 199640 163740 199646
rect 163688 199582 163740 199588
rect 163872 199640 163924 199646
rect 163872 199582 163924 199588
rect 163594 189408 163650 189417
rect 163594 189343 163650 189352
rect 163700 182442 163728 199582
rect 163780 199504 163832 199510
rect 163780 199446 163832 199452
rect 163792 197062 163820 199446
rect 163780 197056 163832 197062
rect 163780 196998 163832 197004
rect 163884 196926 163912 199582
rect 163976 197266 164004 199702
rect 164160 198734 164188 199736
rect 164298 199730 164326 200124
rect 164390 199850 164418 200124
rect 164378 199844 164430 199850
rect 164378 199786 164430 199792
rect 164482 199730 164510 200124
rect 164298 199702 164372 199730
rect 164160 198706 164280 198734
rect 164252 197305 164280 198706
rect 164238 197296 164294 197305
rect 163964 197260 164016 197266
rect 164238 197231 164294 197240
rect 163964 197202 164016 197208
rect 163872 196920 163924 196926
rect 163872 196862 163924 196868
rect 164344 195242 164372 199702
rect 164436 199702 164510 199730
rect 164436 196722 164464 199702
rect 164574 199696 164602 200124
rect 164666 199764 164694 200124
rect 164758 199918 164786 200124
rect 164746 199912 164798 199918
rect 164850 199889 164878 200124
rect 164942 199918 164970 200124
rect 164930 199912 164982 199918
rect 164746 199854 164798 199860
rect 164836 199880 164892 199889
rect 164930 199854 164982 199860
rect 164836 199815 164892 199824
rect 165034 199764 165062 200124
rect 165126 199889 165154 200124
rect 165112 199880 165168 199889
rect 165112 199815 165168 199824
rect 164666 199736 164740 199764
rect 164574 199668 164648 199696
rect 164516 199572 164568 199578
rect 164516 199514 164568 199520
rect 164424 196716 164476 196722
rect 164424 196658 164476 196664
rect 164528 196382 164556 199514
rect 164516 196376 164568 196382
rect 164516 196318 164568 196324
rect 164344 195214 164556 195242
rect 164424 195152 164476 195158
rect 164424 195094 164476 195100
rect 164238 191176 164294 191185
rect 164238 191111 164294 191120
rect 163688 182436 163740 182442
rect 163688 182378 163740 182384
rect 163228 152448 163280 152454
rect 163228 152390 163280 152396
rect 162952 148640 163004 148646
rect 162952 148582 163004 148588
rect 164252 148442 164280 191111
rect 164332 190052 164384 190058
rect 164332 189994 164384 190000
rect 164344 148510 164372 189994
rect 164436 148782 164464 195094
rect 164528 152862 164556 195214
rect 164620 190058 164648 199668
rect 164712 191185 164740 199736
rect 164988 199736 165062 199764
rect 164884 199708 164936 199714
rect 164884 199650 164936 199656
rect 164792 199504 164844 199510
rect 164792 199446 164844 199452
rect 164804 199306 164832 199446
rect 164792 199300 164844 199306
rect 164792 199242 164844 199248
rect 164896 197305 164924 199650
rect 164882 197296 164938 197305
rect 164882 197231 164938 197240
rect 164988 196897 165016 199736
rect 165218 199696 165246 200124
rect 165310 199764 165338 200124
rect 165402 199889 165430 200124
rect 165388 199880 165444 199889
rect 165494 199850 165522 200124
rect 165388 199815 165444 199824
rect 165482 199844 165534 199850
rect 165482 199786 165534 199792
rect 165310 199736 165384 199764
rect 165218 199668 165292 199696
rect 165068 199640 165120 199646
rect 165068 199582 165120 199588
rect 165080 197577 165108 199582
rect 165158 199336 165214 199345
rect 165158 199271 165214 199280
rect 165066 197568 165122 197577
rect 165066 197503 165122 197512
rect 164974 196888 165030 196897
rect 164974 196823 165030 196832
rect 165172 195158 165200 199271
rect 165264 197441 165292 199668
rect 165356 198014 165384 199736
rect 165586 199730 165614 200124
rect 165540 199702 165614 199730
rect 165436 199572 165488 199578
rect 165436 199514 165488 199520
rect 165344 198008 165396 198014
rect 165344 197950 165396 197956
rect 165448 197674 165476 199514
rect 165436 197668 165488 197674
rect 165436 197610 165488 197616
rect 165250 197432 165306 197441
rect 165250 197367 165306 197376
rect 165540 197354 165568 199702
rect 165678 199696 165706 200124
rect 165770 199918 165798 200124
rect 165862 199918 165890 200124
rect 165954 199918 165982 200124
rect 165758 199912 165810 199918
rect 165758 199854 165810 199860
rect 165850 199912 165902 199918
rect 165850 199854 165902 199860
rect 165942 199912 165994 199918
rect 165942 199854 165994 199860
rect 165804 199776 165856 199782
rect 165804 199718 165856 199724
rect 165896 199776 165948 199782
rect 165896 199718 165948 199724
rect 165678 199668 165752 199696
rect 165620 199436 165672 199442
rect 165620 199378 165672 199384
rect 165448 197326 165568 197354
rect 165342 197296 165398 197305
rect 165342 197231 165398 197240
rect 165160 195152 165212 195158
rect 165160 195094 165212 195100
rect 164698 191176 164754 191185
rect 164698 191111 164754 191120
rect 164608 190052 164660 190058
rect 164608 189994 164660 190000
rect 165356 180794 165384 197231
rect 165448 192982 165476 197326
rect 165632 195838 165660 199378
rect 165724 197402 165752 199668
rect 165712 197396 165764 197402
rect 165712 197338 165764 197344
rect 165620 195832 165672 195838
rect 165620 195774 165672 195780
rect 165620 195220 165672 195226
rect 165620 195162 165672 195168
rect 165436 192976 165488 192982
rect 165436 192918 165488 192924
rect 164620 180766 165384 180794
rect 164516 152856 164568 152862
rect 164516 152798 164568 152804
rect 164620 152697 164648 180766
rect 164606 152688 164662 152697
rect 164606 152623 164662 152632
rect 165632 149054 165660 195162
rect 165712 195016 165764 195022
rect 165712 194958 165764 194964
rect 165620 149048 165672 149054
rect 165620 148990 165672 148996
rect 164424 148776 164476 148782
rect 164424 148718 164476 148724
rect 165724 148578 165752 194958
rect 165816 192302 165844 199718
rect 165804 192296 165856 192302
rect 165804 192238 165856 192244
rect 165908 148918 165936 199718
rect 166046 199696 166074 200124
rect 166138 199918 166166 200124
rect 166126 199912 166178 199918
rect 166126 199854 166178 199860
rect 166230 199764 166258 200124
rect 166000 199668 166074 199696
rect 166184 199736 166258 199764
rect 166000 199073 166028 199668
rect 166080 199504 166132 199510
rect 166080 199446 166132 199452
rect 165986 199064 166042 199073
rect 165986 198999 166042 199008
rect 165986 198928 166042 198937
rect 165986 198863 165988 198872
rect 166040 198863 166042 198872
rect 165988 198834 166040 198840
rect 166092 198830 166120 199446
rect 166080 198824 166132 198830
rect 166080 198766 166132 198772
rect 165988 197396 166040 197402
rect 165988 197338 166040 197344
rect 166000 152794 166028 197338
rect 166184 194594 166212 199736
rect 166322 199696 166350 200124
rect 166414 199889 166442 200124
rect 166506 199918 166534 200124
rect 166494 199912 166546 199918
rect 166400 199880 166456 199889
rect 166494 199854 166546 199860
rect 166400 199815 166456 199824
rect 166598 199764 166626 200124
rect 166276 199668 166350 199696
rect 166552 199736 166626 199764
rect 166690 199764 166718 200124
rect 166782 199889 166810 200124
rect 166768 199880 166824 199889
rect 166768 199815 166824 199824
rect 166874 199764 166902 200124
rect 166690 199736 166764 199764
rect 166276 198734 166304 199668
rect 166448 199640 166500 199646
rect 166448 199582 166500 199588
rect 166356 199572 166408 199578
rect 166356 199514 166408 199520
rect 166368 199345 166396 199514
rect 166354 199336 166410 199345
rect 166354 199271 166410 199280
rect 166276 198706 166396 198734
rect 166368 197305 166396 198706
rect 166354 197296 166410 197305
rect 166354 197231 166410 197240
rect 166460 195022 166488 199582
rect 166552 198121 166580 199736
rect 166736 199646 166764 199736
rect 166828 199736 166902 199764
rect 166966 199764 166994 200124
rect 167058 199918 167086 200124
rect 167046 199912 167098 199918
rect 167150 199889 167178 200124
rect 167242 199918 167270 200124
rect 167334 199918 167362 200124
rect 167230 199912 167282 199918
rect 167046 199854 167098 199860
rect 167136 199880 167192 199889
rect 167230 199854 167282 199860
rect 167322 199912 167374 199918
rect 167426 199889 167454 200124
rect 167322 199854 167374 199860
rect 167412 199880 167468 199889
rect 167136 199815 167192 199824
rect 167412 199815 167468 199824
rect 167184 199776 167236 199782
rect 166966 199736 167132 199764
rect 166632 199640 166684 199646
rect 166632 199582 166684 199588
rect 166724 199640 166776 199646
rect 166724 199582 166776 199588
rect 166644 198762 166672 199582
rect 166828 198937 166856 199736
rect 167000 199640 167052 199646
rect 167000 199582 167052 199588
rect 166908 199572 166960 199578
rect 166908 199514 166960 199520
rect 166814 198928 166870 198937
rect 166724 198892 166776 198898
rect 166814 198863 166870 198872
rect 166724 198834 166776 198840
rect 166632 198756 166684 198762
rect 166632 198698 166684 198704
rect 166538 198112 166594 198121
rect 166538 198047 166594 198056
rect 166736 195226 166764 198834
rect 166920 196761 166948 199514
rect 166906 196752 166962 196761
rect 166906 196687 166962 196696
rect 167012 196042 167040 199582
rect 167104 198626 167132 199736
rect 167184 199718 167236 199724
rect 167368 199776 167420 199782
rect 167518 199764 167546 200124
rect 167610 199918 167638 200124
rect 167598 199912 167650 199918
rect 167598 199854 167650 199860
rect 167702 199764 167730 200124
rect 167368 199718 167420 199724
rect 167472 199736 167546 199764
rect 167656 199736 167730 199764
rect 167196 198694 167224 199718
rect 167380 199628 167408 199718
rect 167288 199600 167408 199628
rect 167184 198688 167236 198694
rect 167184 198630 167236 198636
rect 167092 198620 167144 198626
rect 167092 198562 167144 198568
rect 167000 196036 167052 196042
rect 167000 195978 167052 195984
rect 166724 195220 166776 195226
rect 166724 195162 166776 195168
rect 166448 195016 166500 195022
rect 166448 194958 166500 194964
rect 166184 194566 166304 194594
rect 166276 190454 166304 194566
rect 167288 191282 167316 199600
rect 167472 199560 167500 199736
rect 167380 199532 167500 199560
rect 167380 199306 167408 199532
rect 167656 199458 167684 199736
rect 167794 199696 167822 200124
rect 167886 199889 167914 200124
rect 167978 199918 168006 200124
rect 167966 199912 168018 199918
rect 167872 199880 167928 199889
rect 167966 199854 168018 199860
rect 167872 199815 167928 199824
rect 168070 199764 168098 200124
rect 167564 199430 167684 199458
rect 167748 199668 167822 199696
rect 167932 199736 168098 199764
rect 167368 199300 167420 199306
rect 167368 199242 167420 199248
rect 167564 197577 167592 199430
rect 167644 199368 167696 199374
rect 167644 199310 167696 199316
rect 167550 197568 167606 197577
rect 167550 197503 167606 197512
rect 167656 194594 167684 199310
rect 167748 197538 167776 199668
rect 167826 198928 167882 198937
rect 167826 198863 167882 198872
rect 167736 197532 167788 197538
rect 167736 197474 167788 197480
rect 167472 194566 167684 194594
rect 167276 191276 167328 191282
rect 167276 191218 167328 191224
rect 167472 191162 167500 194566
rect 167104 191134 167500 191162
rect 166276 190426 166948 190454
rect 165988 152788 166040 152794
rect 165988 152730 166040 152736
rect 165896 148912 165948 148918
rect 165896 148854 165948 148860
rect 166920 148850 166948 190426
rect 167104 152658 167132 191134
rect 167840 186314 167868 198863
rect 167932 193905 167960 199736
rect 168162 199696 168190 200124
rect 168116 199668 168190 199696
rect 168254 199696 168282 200124
rect 168346 199764 168374 200124
rect 168438 199918 168466 200124
rect 168530 199918 168558 200124
rect 168622 199918 168650 200124
rect 168426 199912 168478 199918
rect 168426 199854 168478 199860
rect 168518 199912 168570 199918
rect 168518 199854 168570 199860
rect 168610 199912 168662 199918
rect 168610 199854 168662 199860
rect 168346 199736 168420 199764
rect 168254 199668 168328 199696
rect 168012 199640 168064 199646
rect 168012 199582 168064 199588
rect 168024 197441 168052 199582
rect 168010 197432 168066 197441
rect 168010 197367 168066 197376
rect 167918 193896 167974 193905
rect 167918 193831 167974 193840
rect 167288 186286 167868 186314
rect 167288 155242 167316 186286
rect 168116 180794 168144 199668
rect 168196 199572 168248 199578
rect 168196 199514 168248 199520
rect 168208 197169 168236 199514
rect 168300 197305 168328 199668
rect 168286 197296 168342 197305
rect 168286 197231 168342 197240
rect 168194 197160 168250 197169
rect 168194 197095 168250 197104
rect 168392 194594 168420 199736
rect 168564 199708 168616 199714
rect 168564 199650 168616 199656
rect 168472 199504 168524 199510
rect 168472 199446 168524 199452
rect 168484 197062 168512 199446
rect 168472 197056 168524 197062
rect 168472 196998 168524 197004
rect 168208 194566 168420 194594
rect 168208 193866 168236 194566
rect 168576 194041 168604 199650
rect 168714 199628 168742 200124
rect 168806 199918 168834 200124
rect 168898 199918 168926 200124
rect 168990 199918 169018 200124
rect 168794 199912 168846 199918
rect 168794 199854 168846 199860
rect 168886 199912 168938 199918
rect 168886 199854 168938 199860
rect 168978 199912 169030 199918
rect 168978 199854 169030 199860
rect 169082 199730 169110 200124
rect 169174 199918 169202 200124
rect 169266 199918 169294 200124
rect 169358 199918 169386 200124
rect 169162 199912 169214 199918
rect 169162 199854 169214 199860
rect 169254 199912 169306 199918
rect 169254 199854 169306 199860
rect 169346 199912 169398 199918
rect 169346 199854 169398 199860
rect 168840 199708 168892 199714
rect 168840 199650 168892 199656
rect 168932 199708 168984 199714
rect 168932 199650 168984 199656
rect 169036 199702 169110 199730
rect 169208 199708 169260 199714
rect 168668 199600 168742 199628
rect 168562 194032 168618 194041
rect 168562 193967 168618 193976
rect 168196 193860 168248 193866
rect 168196 193802 168248 193808
rect 168288 191276 168340 191282
rect 168288 191218 168340 191224
rect 167840 180766 168144 180794
rect 167276 155236 167328 155242
rect 167276 155178 167328 155184
rect 167092 152652 167144 152658
rect 167092 152594 167144 152600
rect 166908 148844 166960 148850
rect 166908 148786 166960 148792
rect 167840 148714 167868 180766
rect 168300 152590 168328 191218
rect 168668 191162 168696 199600
rect 168852 197354 168880 199650
rect 168760 197326 168880 197354
rect 168760 192642 168788 197326
rect 168840 197056 168892 197062
rect 168840 196998 168892 197004
rect 168852 193934 168880 196998
rect 168840 193928 168892 193934
rect 168840 193870 168892 193876
rect 168748 192636 168800 192642
rect 168748 192578 168800 192584
rect 168392 191134 168696 191162
rect 168392 152726 168420 191134
rect 168472 191072 168524 191078
rect 168472 191014 168524 191020
rect 168484 155310 168512 191014
rect 168944 186314 168972 199650
rect 169036 197441 169064 199702
rect 169208 199650 169260 199656
rect 169300 199708 169352 199714
rect 169450 199696 169478 200124
rect 169300 199650 169352 199656
rect 169404 199668 169478 199696
rect 169116 199640 169168 199646
rect 169116 199582 169168 199588
rect 169022 197432 169078 197441
rect 169022 197367 169078 197376
rect 169128 194594 169156 199582
rect 169036 194566 169156 194594
rect 169036 192778 169064 194566
rect 169024 192772 169076 192778
rect 169024 192714 169076 192720
rect 169220 191078 169248 199650
rect 169312 197985 169340 199650
rect 169298 197976 169354 197985
rect 169298 197911 169354 197920
rect 169404 192846 169432 199668
rect 169542 199628 169570 200124
rect 169634 199889 169662 200124
rect 169620 199880 169676 199889
rect 169620 199815 169676 199824
rect 169726 199764 169754 200124
rect 169496 199600 169570 199628
rect 169680 199736 169754 199764
rect 169392 192840 169444 192846
rect 169392 192782 169444 192788
rect 169208 191072 169260 191078
rect 169208 191014 169260 191020
rect 168576 186286 168972 186314
rect 168576 155446 168604 186286
rect 169496 180794 169524 199600
rect 169576 199504 169628 199510
rect 169576 199446 169628 199452
rect 169588 197305 169616 199446
rect 169680 199322 169708 199736
rect 169818 199458 169846 200124
rect 169910 199594 169938 200124
rect 170002 199696 170030 200124
rect 170094 199764 170122 200124
rect 170186 199918 170214 200124
rect 170174 199912 170226 199918
rect 170174 199854 170226 199860
rect 170278 199764 170306 200124
rect 170370 199850 170398 200124
rect 170462 199889 170490 200124
rect 170554 199918 170582 200124
rect 170646 199918 170674 200124
rect 170738 199918 170766 200124
rect 170542 199912 170594 199918
rect 170448 199880 170504 199889
rect 170358 199844 170410 199850
rect 170542 199854 170594 199860
rect 170634 199912 170686 199918
rect 170634 199854 170686 199860
rect 170726 199912 170778 199918
rect 170726 199854 170778 199860
rect 170448 199815 170504 199824
rect 170358 199786 170410 199792
rect 170830 199764 170858 200124
rect 170094 199736 170168 199764
rect 170002 199668 170076 199696
rect 169910 199566 169984 199594
rect 169818 199430 169892 199458
rect 169680 199294 169800 199322
rect 169772 198830 169800 199294
rect 169760 198824 169812 198830
rect 169760 198766 169812 198772
rect 169574 197296 169630 197305
rect 169574 197231 169630 197240
rect 169760 196308 169812 196314
rect 169760 196250 169812 196256
rect 169772 195226 169800 196250
rect 169760 195220 169812 195226
rect 169760 195162 169812 195168
rect 169864 191298 169892 199430
rect 169956 196450 169984 199566
rect 170048 199442 170076 199668
rect 170036 199436 170088 199442
rect 170036 199378 170088 199384
rect 169944 196444 169996 196450
rect 169944 196386 169996 196392
rect 170140 194594 170168 199736
rect 170232 199736 170306 199764
rect 170784 199736 170858 199764
rect 170232 198354 170260 199736
rect 170588 199708 170640 199714
rect 170588 199650 170640 199656
rect 170680 199708 170732 199714
rect 170680 199650 170732 199656
rect 170404 199640 170456 199646
rect 170404 199582 170456 199588
rect 170496 199640 170548 199646
rect 170496 199582 170548 199588
rect 170312 199368 170364 199374
rect 170416 199345 170444 199582
rect 170312 199310 170364 199316
rect 170402 199336 170458 199345
rect 170324 198898 170352 199310
rect 170402 199271 170458 199280
rect 170404 199232 170456 199238
rect 170404 199174 170456 199180
rect 170416 198898 170444 199174
rect 170312 198892 170364 198898
rect 170312 198834 170364 198840
rect 170404 198892 170456 198898
rect 170404 198834 170456 198840
rect 170508 198734 170536 199582
rect 170416 198706 170536 198734
rect 170220 198348 170272 198354
rect 170220 198290 170272 198296
rect 170416 198218 170444 198706
rect 170496 198620 170548 198626
rect 170496 198562 170548 198568
rect 170404 198212 170456 198218
rect 170404 198154 170456 198160
rect 170402 197296 170458 197305
rect 170402 197231 170458 197240
rect 170048 194566 170168 194594
rect 170048 191434 170076 194566
rect 170048 191406 170260 191434
rect 169864 191270 170168 191298
rect 169944 191208 169996 191214
rect 169944 191150 169996 191156
rect 169852 191140 169904 191146
rect 169852 191082 169904 191088
rect 168668 180766 169524 180794
rect 168564 155440 168616 155446
rect 168564 155382 168616 155388
rect 168668 155378 168696 180766
rect 168656 155372 168708 155378
rect 168656 155314 168708 155320
rect 168472 155304 168524 155310
rect 168472 155246 168524 155252
rect 168380 152720 168432 152726
rect 168380 152662 168432 152668
rect 168288 152584 168340 152590
rect 168288 152526 168340 152532
rect 167828 148708 167880 148714
rect 167828 148650 167880 148656
rect 165712 148572 165764 148578
rect 165712 148514 165764 148520
rect 164332 148504 164384 148510
rect 164332 148446 164384 148452
rect 164240 148436 164292 148442
rect 164240 148378 164292 148384
rect 164238 145616 164294 145625
rect 164238 145551 164294 145560
rect 163962 143984 164018 143993
rect 163962 143919 164018 143928
rect 163594 143168 163650 143177
rect 163594 143103 163650 143112
rect 162858 141400 162914 141409
rect 162858 141335 162914 141344
rect 160664 139862 161092 139890
rect 161644 139862 161980 139890
rect 162196 139862 162532 139890
rect 162734 140134 162808 140162
rect 162734 139876 162762 140134
rect 163608 139890 163636 143103
rect 163976 139890 164004 143919
rect 163300 139862 163636 139890
rect 163852 139862 164004 139890
rect 164252 139890 164280 145551
rect 168010 144800 168066 144809
rect 168010 144735 168066 144744
rect 166354 144664 166410 144673
rect 165528 144628 165580 144634
rect 166354 144599 166410 144608
rect 165528 144570 165580 144576
rect 165250 143440 165306 143449
rect 165250 143375 165306 143384
rect 165264 139890 165292 143375
rect 165540 140162 165568 144570
rect 164252 139862 164404 139890
rect 164956 139862 165292 139890
rect 165494 140134 165568 140162
rect 165494 139876 165522 140134
rect 166368 139890 166396 144599
rect 166908 142928 166960 142934
rect 166908 142870 166960 142876
rect 166920 139890 166948 142870
rect 167460 141500 167512 141506
rect 167460 141442 167512 141448
rect 167472 139890 167500 141442
rect 168024 139890 168052 144735
rect 169668 144696 169720 144702
rect 169668 144638 169720 144644
rect 168288 143064 168340 143070
rect 168288 143006 168340 143012
rect 168300 140162 168328 143006
rect 169116 141568 169168 141574
rect 169116 141510 169168 141516
rect 166060 139862 166396 139890
rect 166612 139862 166948 139890
rect 167164 139862 167500 139890
rect 167716 139862 168052 139890
rect 168254 140134 168328 140162
rect 168254 139876 168282 140134
rect 169128 139890 169156 141510
rect 169680 139890 169708 144638
rect 169864 140350 169892 191082
rect 169852 140344 169904 140350
rect 169852 140286 169904 140292
rect 169956 140214 169984 191150
rect 170036 191072 170088 191078
rect 170036 191014 170088 191020
rect 170048 140321 170076 191014
rect 170140 147422 170168 191270
rect 170232 191078 170260 191406
rect 170220 191072 170272 191078
rect 170220 191014 170272 191020
rect 170416 186314 170444 197231
rect 170508 192438 170536 198562
rect 170496 192432 170548 192438
rect 170496 192374 170548 192380
rect 170600 191146 170628 199650
rect 170692 197441 170720 199650
rect 170784 198286 170812 199736
rect 170922 199696 170950 200124
rect 171014 199764 171042 200124
rect 171106 199889 171134 200124
rect 171092 199880 171148 199889
rect 171092 199815 171148 199824
rect 171014 199736 171088 199764
rect 170922 199668 170996 199696
rect 170864 199572 170916 199578
rect 170864 199514 170916 199520
rect 170876 199345 170904 199514
rect 170862 199336 170918 199345
rect 170862 199271 170918 199280
rect 170968 198734 170996 199668
rect 170876 198706 170996 198734
rect 170772 198280 170824 198286
rect 170772 198222 170824 198228
rect 170678 197432 170734 197441
rect 170678 197367 170734 197376
rect 170876 191214 170904 198706
rect 171060 198257 171088 199736
rect 171198 199458 171226 200124
rect 171290 199918 171318 200124
rect 171278 199912 171330 199918
rect 171278 199854 171330 199860
rect 171382 199594 171410 200124
rect 171474 199696 171502 200124
rect 171566 199889 171594 200124
rect 171658 199918 171686 200124
rect 171750 199918 171778 200124
rect 171646 199912 171698 199918
rect 171552 199880 171608 199889
rect 171646 199854 171698 199860
rect 171738 199912 171790 199918
rect 171738 199854 171790 199860
rect 171552 199815 171608 199824
rect 171692 199776 171744 199782
rect 171842 199764 171870 200124
rect 171934 199889 171962 200124
rect 172026 199918 172054 200124
rect 172014 199912 172066 199918
rect 171920 199880 171976 199889
rect 172014 199854 172066 199860
rect 171920 199815 171976 199824
rect 171692 199718 171744 199724
rect 171796 199736 171870 199764
rect 172118 199764 172146 200124
rect 172210 199918 172238 200124
rect 172198 199912 172250 199918
rect 172198 199854 172250 199860
rect 172302 199764 172330 200124
rect 172118 199736 172192 199764
rect 171474 199668 171548 199696
rect 171382 199566 171456 199594
rect 171324 199504 171376 199510
rect 171198 199430 171272 199458
rect 171324 199446 171376 199452
rect 171138 199336 171194 199345
rect 171138 199271 171194 199280
rect 171152 198558 171180 199271
rect 171140 198552 171192 198558
rect 171140 198494 171192 198500
rect 171046 198248 171102 198257
rect 171046 198183 171102 198192
rect 171048 198144 171100 198150
rect 171048 198086 171100 198092
rect 171060 195974 171088 198086
rect 171140 198076 171192 198082
rect 171140 198018 171192 198024
rect 171152 196110 171180 198018
rect 171244 197402 171272 199430
rect 171336 198082 171364 199446
rect 171428 198762 171456 199566
rect 171416 198756 171468 198762
rect 171416 198698 171468 198704
rect 171324 198076 171376 198082
rect 171324 198018 171376 198024
rect 171520 197928 171548 199668
rect 171336 197900 171548 197928
rect 171600 197940 171652 197946
rect 171232 197396 171284 197402
rect 171232 197338 171284 197344
rect 171140 196104 171192 196110
rect 171140 196046 171192 196052
rect 171336 195974 171364 197900
rect 171600 197882 171652 197888
rect 171612 197826 171640 197882
rect 171520 197798 171640 197826
rect 171416 197396 171468 197402
rect 171416 197338 171468 197344
rect 171048 195968 171100 195974
rect 171048 195910 171100 195916
rect 171152 195946 171364 195974
rect 170864 191208 170916 191214
rect 170864 191150 170916 191156
rect 170588 191140 170640 191146
rect 170588 191082 170640 191088
rect 170416 186286 170904 186314
rect 170128 147416 170180 147422
rect 170128 147358 170180 147364
rect 170220 143132 170272 143138
rect 170220 143074 170272 143080
rect 170034 140312 170090 140321
rect 170034 140247 170090 140256
rect 169944 140208 169996 140214
rect 169944 140150 169996 140156
rect 170232 139890 170260 143074
rect 170772 141636 170824 141642
rect 170772 141578 170824 141584
rect 170784 139890 170812 141578
rect 170876 140146 170904 186286
rect 171048 143336 171100 143342
rect 171048 143278 171100 143284
rect 171060 140162 171088 143278
rect 171152 140622 171180 195946
rect 171324 191140 171376 191146
rect 171324 191082 171376 191088
rect 171232 189916 171284 189922
rect 171232 189858 171284 189864
rect 171140 140616 171192 140622
rect 171140 140558 171192 140564
rect 171244 140418 171272 189858
rect 171232 140412 171284 140418
rect 171232 140354 171284 140360
rect 171336 140282 171364 191082
rect 171428 146810 171456 197338
rect 171520 195022 171548 197798
rect 171508 195016 171560 195022
rect 171508 194958 171560 194964
rect 171704 180794 171732 199718
rect 171796 197441 171824 199736
rect 171968 199572 172020 199578
rect 171968 199514 172020 199520
rect 171876 199436 171928 199442
rect 171876 199378 171928 199384
rect 171888 198626 171916 199378
rect 171876 198620 171928 198626
rect 171876 198562 171928 198568
rect 171782 197432 171838 197441
rect 171782 197367 171838 197376
rect 171876 196104 171928 196110
rect 171876 196046 171928 196052
rect 171888 195906 171916 196046
rect 171876 195900 171928 195906
rect 171876 195842 171928 195848
rect 171980 191146 172008 199514
rect 172060 199504 172112 199510
rect 172060 199446 172112 199452
rect 172072 199073 172100 199446
rect 172164 199345 172192 199736
rect 172256 199736 172330 199764
rect 172150 199336 172206 199345
rect 172150 199271 172206 199280
rect 172152 199232 172204 199238
rect 172152 199174 172204 199180
rect 172058 199064 172114 199073
rect 172058 198999 172114 199008
rect 172164 198898 172192 199174
rect 172152 198892 172204 198898
rect 172152 198834 172204 198840
rect 172256 198734 172284 199736
rect 172394 199696 172422 200124
rect 172486 199889 172514 200124
rect 172472 199880 172528 199889
rect 172472 199815 172528 199824
rect 172578 199730 172606 200124
rect 172164 198706 172284 198734
rect 172348 199668 172422 199696
rect 172532 199702 172606 199730
rect 172164 197354 172192 198706
rect 172348 197441 172376 199668
rect 172428 199504 172480 199510
rect 172428 199446 172480 199452
rect 172440 198830 172468 199446
rect 172428 198824 172480 198830
rect 172428 198766 172480 198772
rect 172428 198484 172480 198490
rect 172428 198426 172480 198432
rect 172334 197432 172390 197441
rect 172334 197367 172390 197376
rect 172164 197326 172284 197354
rect 172152 195900 172204 195906
rect 172152 195842 172204 195848
rect 172060 195628 172112 195634
rect 172060 195570 172112 195576
rect 172072 195226 172100 195570
rect 172164 195566 172192 195842
rect 172152 195560 172204 195566
rect 172152 195502 172204 195508
rect 172060 195220 172112 195226
rect 172060 195162 172112 195168
rect 171968 191140 172020 191146
rect 171968 191082 172020 191088
rect 172256 189922 172284 197326
rect 172440 196518 172468 198426
rect 172532 198150 172560 199702
rect 172670 199628 172698 200124
rect 172762 199918 172790 200124
rect 172854 199918 172882 200124
rect 172750 199912 172802 199918
rect 172750 199854 172802 199860
rect 172842 199912 172894 199918
rect 172842 199854 172894 199860
rect 172946 199764 172974 200124
rect 173038 199918 173066 200124
rect 173026 199912 173078 199918
rect 173026 199854 173078 199860
rect 173130 199764 173158 200124
rect 172624 199600 172698 199628
rect 172808 199736 172974 199764
rect 173084 199736 173158 199764
rect 172520 198144 172572 198150
rect 172520 198086 172572 198092
rect 172428 196512 172480 196518
rect 172428 196454 172480 196460
rect 172624 195906 172652 199600
rect 172808 199510 172836 199736
rect 172980 199572 173032 199578
rect 172980 199514 173032 199520
rect 172796 199504 172848 199510
rect 172796 199446 172848 199452
rect 172888 199436 172940 199442
rect 172888 199378 172940 199384
rect 172794 199336 172850 199345
rect 172794 199271 172850 199280
rect 172702 199064 172758 199073
rect 172702 198999 172758 199008
rect 172716 198665 172744 198999
rect 172702 198656 172758 198665
rect 172702 198591 172758 198600
rect 172704 198144 172756 198150
rect 172704 198086 172756 198092
rect 172612 195900 172664 195906
rect 172612 195842 172664 195848
rect 172716 194594 172744 198086
rect 172624 194566 172744 194594
rect 172520 191208 172572 191214
rect 172520 191150 172572 191156
rect 172244 189916 172296 189922
rect 172244 189858 172296 189864
rect 171520 180766 171732 180794
rect 171520 147558 171548 180766
rect 171600 149864 171652 149870
rect 171600 149806 171652 149812
rect 171508 147552 171560 147558
rect 171508 147494 171560 147500
rect 171416 146804 171468 146810
rect 171416 146746 171468 146752
rect 171324 140276 171376 140282
rect 171324 140218 171376 140224
rect 170864 140140 170916 140146
rect 170864 140082 170916 140088
rect 171014 140134 171088 140162
rect 171230 140176 171286 140185
rect 168820 139862 169156 139890
rect 169372 139862 169708 139890
rect 169924 139862 170260 139890
rect 170476 139862 170812 139890
rect 171014 139876 171042 140134
rect 171612 140162 171640 149806
rect 172532 145926 172560 191150
rect 172624 147150 172652 194566
rect 172704 191140 172756 191146
rect 172704 191082 172756 191088
rect 172716 147257 172744 191082
rect 172702 147248 172758 147257
rect 172702 147183 172758 147192
rect 172612 147144 172664 147150
rect 172612 147086 172664 147092
rect 172808 146878 172836 199271
rect 172900 197849 172928 199378
rect 172992 199345 173020 199514
rect 172978 199336 173034 199345
rect 172978 199271 173034 199280
rect 172980 198824 173032 198830
rect 172980 198766 173032 198772
rect 172886 197840 172942 197849
rect 172886 197775 172942 197784
rect 172992 197305 173020 198766
rect 172978 197296 173034 197305
rect 172978 197231 173034 197240
rect 172888 195900 172940 195906
rect 172888 195842 172940 195848
rect 172900 192914 172928 195842
rect 172888 192908 172940 192914
rect 172888 192850 172940 192856
rect 173084 180794 173112 199736
rect 173222 199696 173250 200124
rect 173314 199918 173342 200124
rect 173302 199912 173354 199918
rect 173302 199854 173354 199860
rect 173406 199764 173434 200124
rect 173176 199668 173250 199696
rect 173360 199736 173434 199764
rect 173498 199764 173526 200124
rect 173590 199918 173618 200124
rect 173578 199912 173630 199918
rect 173578 199854 173630 199860
rect 173682 199764 173710 200124
rect 173774 199889 173802 200124
rect 173866 199918 173894 200124
rect 173958 199918 173986 200124
rect 173854 199912 173906 199918
rect 173760 199880 173816 199889
rect 173854 199854 173906 199860
rect 173946 199912 173998 199918
rect 173946 199854 173998 199860
rect 173760 199815 173816 199824
rect 173498 199736 173572 199764
rect 173176 197305 173204 199668
rect 173256 198824 173308 198830
rect 173254 198792 173256 198801
rect 173308 198792 173310 198801
rect 173254 198727 173310 198736
rect 173256 198076 173308 198082
rect 173256 198018 173308 198024
rect 173162 197296 173218 197305
rect 173162 197231 173218 197240
rect 173268 194594 173296 198018
rect 173176 194566 173296 194594
rect 173176 192681 173204 194566
rect 173162 192672 173218 192681
rect 173162 192607 173218 192616
rect 173360 191214 173388 199736
rect 173440 199504 173492 199510
rect 173440 199446 173492 199452
rect 173452 198529 173480 199446
rect 173438 198520 173494 198529
rect 173438 198455 173494 198464
rect 173440 198416 173492 198422
rect 173440 198358 173492 198364
rect 173452 196450 173480 198358
rect 173544 197441 173572 199736
rect 173636 199736 173710 199764
rect 173530 197432 173586 197441
rect 173530 197367 173586 197376
rect 173440 196444 173492 196450
rect 173440 196386 173492 196392
rect 173348 191208 173400 191214
rect 173348 191150 173400 191156
rect 173636 191146 173664 199736
rect 174050 199730 174078 200124
rect 174142 199850 174170 200124
rect 174234 199889 174262 200124
rect 174220 199880 174276 199889
rect 174130 199844 174182 199850
rect 174220 199815 174276 199824
rect 174130 199786 174182 199792
rect 174050 199702 174124 199730
rect 173992 199640 174044 199646
rect 173992 199582 174044 199588
rect 173808 199572 173860 199578
rect 173808 199514 173860 199520
rect 173900 199572 173952 199578
rect 173900 199514 173952 199520
rect 173716 199504 173768 199510
rect 173716 199446 173768 199452
rect 173728 197985 173756 199446
rect 173714 197976 173770 197985
rect 173714 197911 173770 197920
rect 173820 197878 173848 199514
rect 173912 198150 173940 199514
rect 173900 198144 173952 198150
rect 173900 198086 173952 198092
rect 173808 197872 173860 197878
rect 173808 197814 173860 197820
rect 173716 197804 173768 197810
rect 173716 197746 173768 197752
rect 173728 195906 173756 197746
rect 173716 195900 173768 195906
rect 173716 195842 173768 195848
rect 174004 194594 174032 199582
rect 174096 197402 174124 199702
rect 174176 199640 174228 199646
rect 174326 199628 174354 200124
rect 174418 199696 174446 200124
rect 174510 199764 174538 200124
rect 174602 199918 174630 200124
rect 174694 199918 174722 200124
rect 174590 199912 174642 199918
rect 174590 199854 174642 199860
rect 174682 199912 174734 199918
rect 174682 199854 174734 199860
rect 174786 199764 174814 200124
rect 174510 199736 174584 199764
rect 174418 199668 174492 199696
rect 174326 199600 174400 199628
rect 174176 199582 174228 199588
rect 174188 198801 174216 199582
rect 174266 199472 174322 199481
rect 174266 199407 174322 199416
rect 174174 198792 174230 198801
rect 174174 198727 174230 198736
rect 174176 198688 174228 198694
rect 174176 198630 174228 198636
rect 174188 198490 174216 198630
rect 174176 198484 174228 198490
rect 174176 198426 174228 198432
rect 174176 198008 174228 198014
rect 174176 197950 174228 197956
rect 174084 197396 174136 197402
rect 174084 197338 174136 197344
rect 174188 196790 174216 197950
rect 174176 196784 174228 196790
rect 174176 196726 174228 196732
rect 174004 194566 174216 194594
rect 174084 191208 174136 191214
rect 174084 191150 174136 191156
rect 173624 191140 173676 191146
rect 173624 191082 173676 191088
rect 173992 191140 174044 191146
rect 173992 191082 174044 191088
rect 173900 191072 173952 191078
rect 173900 191014 173952 191020
rect 172900 180766 173112 180794
rect 172900 147082 172928 180766
rect 172980 147212 173032 147218
rect 172980 147154 173032 147160
rect 172888 147076 172940 147082
rect 172888 147018 172940 147024
rect 172796 146872 172848 146878
rect 172796 146814 172848 146820
rect 172520 145920 172572 145926
rect 172520 145862 172572 145868
rect 172428 144832 172480 144838
rect 172428 144774 172480 144780
rect 171230 140111 171286 140120
rect 171566 140134 171640 140162
rect 171244 139777 171272 140111
rect 171566 139876 171594 140134
rect 172440 139890 172468 144774
rect 172888 143404 172940 143410
rect 172888 143346 172940 143352
rect 172900 139890 172928 143346
rect 172132 139862 172468 139890
rect 172684 139862 172928 139890
rect 172992 139890 173020 147154
rect 173808 144764 173860 144770
rect 173808 144706 173860 144712
rect 173820 140162 173848 144706
rect 173912 140690 173940 191014
rect 174004 145858 174032 191082
rect 174096 146169 174124 191150
rect 174188 147665 174216 194566
rect 174280 186314 174308 199407
rect 174372 197577 174400 199600
rect 174464 199073 174492 199668
rect 174450 199064 174506 199073
rect 174450 198999 174506 199008
rect 174452 198892 174504 198898
rect 174452 198834 174504 198840
rect 174464 198354 174492 198834
rect 174452 198348 174504 198354
rect 174452 198290 174504 198296
rect 174358 197568 174414 197577
rect 174358 197503 174414 197512
rect 174360 197396 174412 197402
rect 174360 197338 174412 197344
rect 174372 192545 174400 197338
rect 174556 194594 174584 199736
rect 174740 199736 174814 199764
rect 174878 199764 174906 200124
rect 174970 199918 174998 200124
rect 174958 199912 175010 199918
rect 175062 199889 175090 200124
rect 175154 199918 175182 200124
rect 175142 199912 175194 199918
rect 174958 199854 175010 199860
rect 175048 199880 175104 199889
rect 175142 199854 175194 199860
rect 175048 199815 175104 199824
rect 175246 199764 175274 200124
rect 175338 199918 175366 200124
rect 175326 199912 175378 199918
rect 175326 199854 175378 199860
rect 175430 199764 175458 200124
rect 175522 199918 175550 200124
rect 175510 199912 175562 199918
rect 175614 199889 175642 200124
rect 175510 199854 175562 199860
rect 175600 199880 175656 199889
rect 175600 199815 175656 199824
rect 175706 199764 175734 200124
rect 174878 199736 174952 199764
rect 174636 199708 174688 199714
rect 174636 199650 174688 199656
rect 174648 198830 174676 199650
rect 174636 198824 174688 198830
rect 174636 198766 174688 198772
rect 174464 194566 174584 194594
rect 174358 192536 174414 192545
rect 174358 192471 174414 192480
rect 174464 191146 174492 194566
rect 174740 191214 174768 199736
rect 174820 199640 174872 199646
rect 174820 199582 174872 199588
rect 174832 199481 174860 199582
rect 174818 199472 174874 199481
rect 174818 199407 174874 199416
rect 174820 198892 174872 198898
rect 174820 198834 174872 198840
rect 174832 198393 174860 198834
rect 174818 198384 174874 198393
rect 174818 198319 174874 198328
rect 174924 197441 174952 199736
rect 175200 199736 175274 199764
rect 175384 199736 175458 199764
rect 175568 199736 175734 199764
rect 175096 199572 175148 199578
rect 175096 199514 175148 199520
rect 175004 199504 175056 199510
rect 175004 199446 175056 199452
rect 175016 197985 175044 199446
rect 175002 197976 175058 197985
rect 175002 197911 175058 197920
rect 174910 197432 174966 197441
rect 174910 197367 174966 197376
rect 175002 197296 175058 197305
rect 175002 197231 175058 197240
rect 174728 191208 174780 191214
rect 174728 191150 174780 191156
rect 174452 191140 174504 191146
rect 174452 191082 174504 191088
rect 175016 191078 175044 197231
rect 175108 195809 175136 199514
rect 175094 195800 175150 195809
rect 175094 195735 175150 195744
rect 175200 195265 175228 199736
rect 175280 199640 175332 199646
rect 175280 199582 175332 199588
rect 175292 197606 175320 199582
rect 175280 197600 175332 197606
rect 175280 197542 175332 197548
rect 175280 197396 175332 197402
rect 175280 197338 175332 197344
rect 175186 195256 175242 195265
rect 175186 195191 175242 195200
rect 175004 191072 175056 191078
rect 175004 191014 175056 191020
rect 174280 186286 174400 186314
rect 174174 147656 174230 147665
rect 174174 147591 174230 147600
rect 174372 147529 174400 186286
rect 174358 147520 174414 147529
rect 174358 147455 174414 147464
rect 174082 146160 174138 146169
rect 174082 146095 174138 146104
rect 175292 145994 175320 197338
rect 175384 197334 175412 199736
rect 175462 199064 175518 199073
rect 175462 198999 175518 199008
rect 175476 198898 175504 198999
rect 175464 198892 175516 198898
rect 175464 198834 175516 198840
rect 175568 198734 175596 199736
rect 175798 199696 175826 200124
rect 175660 199668 175826 199696
rect 175660 198914 175688 199668
rect 175890 199560 175918 200124
rect 175982 199764 176010 200124
rect 176074 199918 176102 200124
rect 176062 199912 176114 199918
rect 176062 199854 176114 199860
rect 175982 199736 176056 199764
rect 175844 199532 175918 199560
rect 175660 198886 175780 198914
rect 175752 198830 175780 198886
rect 175648 198824 175700 198830
rect 175648 198766 175700 198772
rect 175740 198824 175792 198830
rect 175740 198766 175792 198772
rect 175476 198706 175596 198734
rect 175372 197328 175424 197334
rect 175476 197305 175504 198706
rect 175660 198014 175688 198766
rect 175648 198008 175700 198014
rect 175648 197950 175700 197956
rect 175556 197600 175608 197606
rect 175556 197542 175608 197548
rect 175372 197270 175424 197276
rect 175462 197296 175518 197305
rect 175462 197231 175518 197240
rect 175568 197180 175596 197542
rect 175844 197402 175872 199532
rect 175924 198756 175976 198762
rect 175924 198698 175976 198704
rect 175832 197396 175884 197402
rect 175832 197338 175884 197344
rect 175476 197152 175596 197180
rect 175372 191140 175424 191146
rect 175372 191082 175424 191088
rect 175384 146033 175412 191082
rect 175476 149938 175504 197152
rect 175936 194594 175964 198698
rect 176028 197441 176056 199736
rect 176166 199730 176194 200124
rect 176258 199918 176286 200124
rect 176246 199912 176298 199918
rect 176246 199854 176298 199860
rect 176120 199702 176194 199730
rect 176014 197432 176070 197441
rect 176014 197367 176070 197376
rect 175568 194566 175964 194594
rect 175464 149932 175516 149938
rect 175464 149874 175516 149880
rect 175370 146024 175426 146033
rect 175280 145988 175332 145994
rect 175370 145959 175426 145968
rect 175280 145930 175332 145936
rect 175568 145897 175596 194566
rect 176120 191146 176148 199702
rect 176200 199640 176252 199646
rect 176200 199582 176252 199588
rect 176212 199073 176240 199582
rect 176350 199492 176378 200124
rect 176442 199918 176470 200124
rect 176430 199912 176482 199918
rect 176430 199854 176482 199860
rect 176534 199764 176562 200124
rect 176626 199889 176654 200124
rect 176718 199918 176746 200124
rect 176706 199912 176758 199918
rect 176612 199880 176668 199889
rect 176810 199889 176838 200124
rect 176902 199918 176930 200124
rect 176994 199918 177022 200124
rect 177086 199918 177114 200124
rect 176890 199912 176942 199918
rect 176706 199854 176758 199860
rect 176796 199880 176852 199889
rect 176612 199815 176668 199824
rect 176890 199854 176942 199860
rect 176982 199912 177034 199918
rect 176982 199854 177034 199860
rect 177074 199912 177126 199918
rect 177074 199854 177126 199860
rect 176796 199815 176852 199824
rect 177028 199776 177080 199782
rect 176534 199736 176608 199764
rect 176476 199640 176528 199646
rect 176476 199582 176528 199588
rect 176304 199464 176378 199492
rect 176198 199064 176254 199073
rect 176198 198999 176254 199008
rect 176304 195673 176332 199464
rect 176488 199424 176516 199582
rect 176396 199396 176516 199424
rect 176290 195664 176346 195673
rect 176290 195599 176346 195608
rect 176108 191140 176160 191146
rect 176108 191082 176160 191088
rect 176396 180794 176424 199396
rect 176474 199064 176530 199073
rect 176474 198999 176530 199008
rect 176488 198762 176516 198999
rect 176476 198756 176528 198762
rect 176476 198698 176528 198704
rect 176580 198529 176608 199736
rect 177178 199764 177206 200124
rect 177028 199718 177080 199724
rect 177132 199736 177206 199764
rect 176660 199708 176712 199714
rect 176660 199650 176712 199656
rect 176936 199708 176988 199714
rect 176936 199650 176988 199656
rect 176566 198520 176622 198529
rect 176566 198455 176622 198464
rect 176672 197334 176700 199650
rect 176844 199572 176896 199578
rect 176844 199514 176896 199520
rect 176752 198824 176804 198830
rect 176752 198766 176804 198772
rect 176568 197328 176620 197334
rect 176568 197270 176620 197276
rect 176660 197328 176712 197334
rect 176660 197270 176712 197276
rect 176580 192817 176608 197270
rect 176764 197169 176792 198766
rect 176750 197160 176806 197169
rect 176750 197095 176806 197104
rect 176856 195945 176884 199514
rect 176842 195936 176898 195945
rect 176842 195871 176898 195880
rect 176844 195220 176896 195226
rect 176844 195162 176896 195168
rect 176752 195152 176804 195158
rect 176752 195094 176804 195100
rect 176660 195084 176712 195090
rect 176660 195026 176712 195032
rect 176566 192808 176622 192817
rect 176566 192743 176622 192752
rect 175660 180766 176424 180794
rect 175660 150006 175688 180766
rect 175648 150000 175700 150006
rect 175648 149942 175700 149948
rect 175554 145888 175610 145897
rect 173992 145852 174044 145858
rect 175554 145823 175610 145832
rect 173992 145794 174044 145800
rect 176292 143472 176344 143478
rect 176292 143414 176344 143420
rect 175740 143268 175792 143274
rect 175740 143210 175792 143216
rect 174636 142996 174688 143002
rect 174636 142938 174688 142944
rect 173900 140684 173952 140690
rect 173900 140626 173952 140632
rect 173774 140134 173848 140162
rect 172992 139862 173236 139890
rect 173774 139876 173802 140134
rect 174648 139890 174676 142938
rect 175188 141704 175240 141710
rect 175188 141646 175240 141652
rect 175200 139890 175228 141646
rect 175752 139890 175780 143210
rect 176304 139890 176332 143414
rect 176568 143200 176620 143206
rect 176568 143142 176620 143148
rect 176580 140162 176608 143142
rect 176672 141273 176700 195026
rect 176658 141264 176714 141273
rect 176658 141199 176714 141208
rect 176764 141137 176792 195094
rect 176856 150142 176884 195162
rect 176844 150136 176896 150142
rect 176844 150078 176896 150084
rect 176948 150074 176976 199650
rect 177040 192953 177068 199718
rect 177132 195129 177160 199736
rect 177270 199696 177298 200124
rect 177224 199668 177298 199696
rect 177362 199696 177390 200124
rect 177454 199764 177482 200124
rect 177546 199866 177574 200124
rect 177652 200110 177804 200138
rect 177546 199838 177620 199866
rect 177454 199736 177528 199764
rect 177362 199668 177436 199696
rect 177224 195226 177252 199668
rect 177304 199572 177356 199578
rect 177304 199514 177356 199520
rect 177316 199345 177344 199514
rect 177302 199336 177358 199345
rect 177302 199271 177358 199280
rect 177408 198121 177436 199668
rect 177394 198112 177450 198121
rect 177394 198047 177450 198056
rect 177500 197985 177528 199736
rect 177486 197976 177542 197985
rect 177486 197911 177542 197920
rect 177304 195560 177356 195566
rect 177304 195502 177356 195508
rect 177316 195226 177344 195502
rect 177212 195220 177264 195226
rect 177212 195162 177264 195168
rect 177304 195220 177356 195226
rect 177304 195162 177356 195168
rect 177592 195158 177620 199838
rect 177672 199504 177724 199510
rect 177672 199446 177724 199452
rect 177684 198762 177712 199446
rect 177672 198756 177724 198762
rect 177672 198698 177724 198704
rect 177776 198098 177804 200110
rect 178314 200087 178370 200096
rect 178500 200116 178552 200122
rect 178132 200048 178184 200054
rect 178132 199990 178184 199996
rect 177948 199980 178000 199986
rect 177948 199922 178000 199928
rect 177854 199880 177910 199889
rect 177854 199815 177910 199824
rect 177684 198070 177804 198098
rect 177580 195152 177632 195158
rect 177118 195120 177174 195129
rect 177580 195094 177632 195100
rect 177684 195090 177712 198070
rect 177118 195055 177174 195064
rect 177672 195084 177724 195090
rect 177672 195026 177724 195032
rect 177868 194594 177896 199815
rect 177960 198830 177988 199922
rect 177948 198824 178000 198830
rect 177948 198766 178000 198772
rect 178144 198529 178172 199990
rect 178130 198520 178186 198529
rect 178328 198490 178356 200087
rect 178500 200058 178552 200064
rect 178130 198455 178186 198464
rect 178316 198484 178368 198490
rect 178316 198426 178368 198432
rect 178512 198014 178540 200058
rect 178500 198008 178552 198014
rect 178500 197950 178552 197956
rect 177776 194566 177896 194594
rect 177776 193089 177804 194566
rect 177762 193080 177818 193089
rect 177762 193015 177818 193024
rect 177026 192944 177082 192953
rect 177026 192879 177082 192888
rect 176936 150068 176988 150074
rect 176936 150010 176988 150016
rect 178408 147484 178460 147490
rect 178408 147426 178460 147432
rect 178224 147348 178276 147354
rect 178224 147290 178276 147296
rect 178040 146736 178092 146742
rect 178040 146678 178092 146684
rect 178052 143426 178080 146678
rect 177960 143398 178080 143426
rect 177396 142724 177448 142730
rect 177396 142666 177448 142672
rect 176750 141128 176806 141137
rect 176750 141063 176806 141072
rect 174340 139862 174676 139890
rect 174892 139862 175228 139890
rect 175444 139862 175780 139890
rect 175996 139862 176332 139890
rect 176534 140134 176608 140162
rect 176534 139876 176562 140134
rect 177408 139890 177436 142666
rect 177960 139890 177988 143398
rect 178236 143018 178264 147290
rect 178316 146124 178368 146130
rect 178316 146066 178368 146072
rect 178052 142990 178264 143018
rect 178052 140758 178080 142990
rect 178132 142792 178184 142798
rect 178132 142734 178184 142740
rect 178040 140752 178092 140758
rect 178040 140694 178092 140700
rect 178144 140554 178172 142734
rect 178224 142588 178276 142594
rect 178224 142530 178276 142536
rect 178236 142225 178264 142530
rect 178222 142216 178278 142225
rect 178222 142151 178278 142160
rect 178132 140548 178184 140554
rect 178132 140490 178184 140496
rect 178038 140176 178094 140185
rect 178038 140111 178094 140120
rect 177100 139862 177436 139890
rect 177652 139862 177988 139890
rect 171230 139768 171286 139777
rect 171230 139703 171286 139712
rect 178052 139602 178080 140111
rect 178328 139754 178356 146066
rect 178420 143342 178448 147426
rect 178696 147286 178724 200631
rect 178684 147280 178736 147286
rect 178684 147222 178736 147228
rect 178788 147218 178816 200670
rect 178960 200456 179012 200462
rect 178960 200398 179012 200404
rect 180248 200456 180300 200462
rect 180248 200398 180300 200404
rect 178972 198734 179000 200398
rect 179328 199436 179380 199442
rect 179328 199378 179380 199384
rect 178880 198706 179000 198734
rect 178776 147212 178828 147218
rect 178776 147154 178828 147160
rect 178880 147098 178908 198706
rect 179340 197946 179368 199378
rect 180156 199232 180208 199238
rect 180156 199174 180208 199180
rect 179328 197940 179380 197946
rect 179328 197882 179380 197888
rect 179052 197736 179104 197742
rect 179052 197678 179104 197684
rect 178960 197668 179012 197674
rect 178960 197610 179012 197616
rect 178972 197062 179000 197610
rect 178960 197056 179012 197062
rect 178960 196998 179012 197004
rect 178960 192296 179012 192302
rect 178960 192238 179012 192244
rect 178512 147070 178908 147098
rect 178408 143336 178460 143342
rect 178408 143278 178460 143284
rect 178512 140434 178540 147070
rect 178868 147008 178920 147014
rect 178868 146950 178920 146956
rect 178592 146056 178644 146062
rect 178592 145998 178644 146004
rect 178604 142798 178632 145998
rect 178592 142792 178644 142798
rect 178592 142734 178644 142740
rect 178592 140548 178644 140554
rect 178592 140490 178644 140496
rect 178204 139726 178356 139754
rect 178420 140406 178540 140434
rect 178040 139596 178092 139602
rect 178040 139538 178092 139544
rect 178420 139369 178448 140406
rect 178604 139890 178632 140490
rect 178604 139862 178756 139890
rect 178880 139369 178908 146950
rect 178972 142154 179000 192238
rect 179064 147014 179092 197678
rect 179144 197328 179196 197334
rect 179144 197270 179196 197276
rect 179156 150385 179184 197270
rect 179694 193216 179750 193225
rect 179236 193180 179288 193186
rect 179694 193151 179750 193160
rect 179236 193122 179288 193128
rect 179142 150376 179198 150385
rect 179142 150311 179198 150320
rect 179248 148306 179276 193122
rect 179708 192710 179736 193151
rect 179696 192704 179748 192710
rect 179696 192646 179748 192652
rect 180064 186924 180116 186930
rect 180064 186866 180116 186872
rect 179236 148300 179288 148306
rect 179236 148242 179288 148248
rect 179144 147620 179196 147626
rect 179144 147562 179196 147568
rect 179052 147008 179104 147014
rect 179052 146950 179104 146956
rect 179156 143478 179184 147562
rect 179236 147552 179288 147558
rect 179236 147494 179288 147500
rect 179328 147552 179380 147558
rect 179328 147494 179380 147500
rect 179248 147286 179276 147494
rect 179236 147280 179288 147286
rect 179236 147222 179288 147228
rect 179236 147144 179288 147150
rect 179236 147086 179288 147092
rect 179248 146810 179276 147086
rect 179236 146804 179288 146810
rect 179236 146746 179288 146752
rect 179144 143472 179196 143478
rect 179144 143414 179196 143420
rect 179340 143410 179368 147494
rect 179512 146260 179564 146266
rect 179512 146202 179564 146208
rect 179420 145512 179472 145518
rect 179420 145454 179472 145460
rect 179328 143404 179380 143410
rect 179328 143346 179380 143352
rect 179432 143274 179460 145454
rect 179420 143268 179472 143274
rect 179420 143210 179472 143216
rect 179524 142730 179552 146202
rect 179604 145444 179656 145450
rect 179604 145386 179656 145392
rect 179512 142724 179564 142730
rect 179512 142666 179564 142672
rect 179616 142154 179644 145386
rect 180076 142154 180104 186866
rect 178972 142126 179092 142154
rect 178960 140752 179012 140758
rect 178960 140694 179012 140700
rect 178972 139890 179000 140694
rect 179064 140486 179092 142126
rect 179432 142126 179644 142154
rect 179984 142126 180104 142154
rect 179144 140684 179196 140690
rect 179144 140626 179196 140632
rect 179052 140480 179104 140486
rect 179052 140422 179104 140428
rect 179156 140049 179184 140626
rect 179142 140040 179198 140049
rect 179142 139975 179198 139984
rect 179432 139890 179460 142126
rect 179512 141772 179564 141778
rect 179512 141714 179564 141720
rect 179524 141098 179552 141714
rect 179512 141092 179564 141098
rect 179512 141034 179564 141040
rect 179984 140554 180012 142126
rect 180168 141545 180196 199174
rect 180260 195974 180288 200398
rect 186780 200184 186832 200190
rect 186780 200126 186832 200132
rect 182916 199504 182968 199510
rect 182916 199446 182968 199452
rect 180892 199436 180944 199442
rect 180892 199378 180944 199384
rect 180800 199232 180852 199238
rect 180800 199174 180852 199180
rect 180812 198898 180840 199174
rect 180800 198892 180852 198898
rect 180800 198834 180852 198840
rect 180616 197532 180668 197538
rect 180616 197474 180668 197480
rect 180524 196376 180576 196382
rect 180524 196318 180576 196324
rect 180260 195946 180380 195974
rect 180248 195696 180300 195702
rect 180248 195638 180300 195644
rect 180154 141536 180210 141545
rect 180154 141471 180210 141480
rect 179972 140548 180024 140554
rect 179972 140490 180024 140496
rect 178972 139862 179308 139890
rect 179432 139862 179860 139890
rect 180260 139369 180288 195638
rect 180352 144158 180380 195946
rect 180432 194948 180484 194954
rect 180432 194890 180484 194896
rect 180340 144152 180392 144158
rect 180340 144094 180392 144100
rect 180444 143478 180472 194890
rect 180536 146878 180564 196318
rect 180628 192370 180656 197474
rect 180904 195974 180932 199378
rect 182824 196240 182876 196246
rect 182824 196182 182876 196188
rect 180812 195946 180932 195974
rect 180616 192364 180668 192370
rect 180616 192306 180668 192312
rect 180524 146872 180576 146878
rect 180524 146814 180576 146820
rect 180432 143472 180484 143478
rect 180432 143414 180484 143420
rect 180340 141772 180392 141778
rect 180340 141714 180392 141720
rect 180352 139890 180380 141714
rect 180812 140729 180840 195946
rect 181536 193112 181588 193118
rect 181536 193054 181588 193060
rect 180892 148368 180944 148374
rect 180892 148310 180944 148316
rect 180798 140720 180854 140729
rect 180798 140655 180854 140664
rect 180904 139890 180932 148310
rect 181548 143342 181576 193054
rect 181628 193044 181680 193050
rect 181628 192986 181680 192992
rect 181536 143336 181588 143342
rect 181536 143278 181588 143284
rect 181166 140720 181222 140729
rect 181166 140655 181222 140664
rect 181180 139890 181208 140655
rect 180352 139862 180412 139890
rect 180904 139862 180964 139890
rect 181180 139862 181516 139890
rect 181272 139505 181300 139862
rect 181640 139602 181668 192986
rect 182272 144968 182324 144974
rect 182272 144910 182324 144916
rect 181996 141840 182048 141846
rect 181996 141782 182048 141788
rect 181810 139904 181866 139913
rect 181810 139839 181866 139848
rect 181628 139596 181680 139602
rect 181628 139538 181680 139544
rect 181824 139534 181852 139839
rect 181902 139768 181958 139777
rect 182008 139754 182036 141782
rect 182284 139890 182312 144910
rect 182284 139862 182620 139890
rect 181958 139726 182068 139754
rect 181902 139703 181958 139712
rect 181902 139632 181958 139641
rect 181902 139567 181958 139576
rect 181812 139528 181864 139534
rect 181258 139496 181314 139505
rect 181812 139470 181864 139476
rect 181916 139466 181944 139567
rect 182836 139505 182864 196182
rect 182928 140962 182956 199446
rect 183836 198824 183888 198830
rect 183836 198766 183888 198772
rect 183192 196172 183244 196178
rect 183192 196114 183244 196120
rect 183008 195764 183060 195770
rect 183008 195706 183060 195712
rect 182916 140956 182968 140962
rect 182916 140898 182968 140904
rect 182928 139890 182956 140898
rect 183020 140010 183048 195706
rect 183204 141914 183232 196114
rect 183284 195832 183336 195838
rect 183284 195774 183336 195780
rect 183192 141908 183244 141914
rect 183192 141850 183244 141856
rect 183008 140004 183060 140010
rect 183008 139946 183060 139952
rect 182928 139862 183172 139890
rect 182822 139496 182878 139505
rect 181258 139431 181314 139440
rect 181904 139460 181956 139466
rect 183296 139466 183324 195774
rect 183848 151814 183876 198766
rect 186688 197940 186740 197946
rect 186688 197882 186740 197888
rect 186596 195288 186648 195294
rect 186596 195230 186648 195236
rect 184664 153196 184716 153202
rect 184664 153138 184716 153144
rect 184204 153128 184256 153134
rect 184204 153070 184256 153076
rect 183848 151786 183968 151814
rect 183836 146192 183888 146198
rect 183836 146134 183888 146140
rect 183468 145580 183520 145586
rect 183468 145522 183520 145528
rect 183480 144974 183508 145522
rect 183468 144968 183520 144974
rect 183848 144945 183876 146134
rect 183468 144910 183520 144916
rect 183834 144936 183890 144945
rect 183834 144871 183890 144880
rect 183744 143268 183796 143274
rect 183744 143210 183796 143216
rect 183756 142186 183784 143210
rect 183744 142180 183796 142186
rect 183744 142122 183796 142128
rect 183756 140162 183784 142122
rect 183710 140134 183784 140162
rect 183710 139876 183738 140134
rect 183848 139890 183876 144871
rect 183940 140729 183968 151786
rect 184112 143064 184164 143070
rect 184112 143006 184164 143012
rect 184124 142798 184152 143006
rect 184112 142792 184164 142798
rect 184112 142734 184164 142740
rect 184216 141982 184244 153070
rect 184296 152448 184348 152454
rect 184296 152390 184348 152396
rect 184308 143070 184336 152390
rect 184388 150340 184440 150346
rect 184388 150282 184440 150288
rect 184296 143064 184348 143070
rect 184296 143006 184348 143012
rect 184204 141976 184256 141982
rect 184204 141918 184256 141924
rect 183926 140720 183982 140729
rect 183926 140655 183982 140664
rect 184400 140457 184428 150282
rect 184572 150272 184624 150278
rect 184572 150214 184624 150220
rect 184480 149660 184532 149666
rect 184480 149602 184532 149608
rect 184492 140622 184520 149602
rect 184480 140616 184532 140622
rect 184480 140558 184532 140564
rect 184386 140448 184442 140457
rect 184386 140383 184442 140392
rect 184584 139942 184612 150214
rect 184676 144906 184704 153138
rect 185584 153060 185636 153066
rect 185584 153002 185636 153008
rect 184756 150204 184808 150210
rect 184756 150146 184808 150152
rect 184664 144900 184716 144906
rect 184664 144842 184716 144848
rect 184768 141166 184796 150146
rect 185030 143304 185086 143313
rect 185030 143239 185086 143248
rect 185044 142769 185072 143239
rect 185030 142760 185086 142769
rect 185030 142695 185086 142704
rect 185032 141228 185084 141234
rect 185032 141170 185084 141176
rect 184756 141160 184808 141166
rect 184756 141102 184808 141108
rect 185044 141030 185072 141170
rect 185596 141114 185624 153002
rect 185768 152992 185820 152998
rect 185768 152934 185820 152940
rect 185780 151814 185808 152934
rect 185780 151786 185900 151814
rect 185768 150408 185820 150414
rect 185768 150350 185820 150356
rect 185676 143404 185728 143410
rect 185676 143346 185728 143352
rect 185688 141234 185716 143346
rect 185676 141228 185728 141234
rect 185676 141170 185728 141176
rect 185596 141086 185716 141114
rect 185032 141024 185084 141030
rect 185032 140966 185084 140972
rect 184754 140720 184810 140729
rect 184754 140655 184810 140664
rect 184664 140072 184716 140078
rect 184664 140014 184716 140020
rect 184572 139936 184624 139942
rect 183848 139862 184276 139890
rect 184572 139878 184624 139884
rect 184676 139505 184704 140014
rect 184768 139890 184796 140655
rect 185044 139890 185072 140966
rect 185584 140208 185636 140214
rect 185584 140150 185636 140156
rect 184768 139862 184828 139890
rect 185044 139862 185380 139890
rect 185596 139874 185624 140150
rect 185688 140078 185716 141086
rect 185676 140072 185728 140078
rect 185676 140014 185728 140020
rect 185584 139868 185636 139874
rect 185584 139810 185636 139816
rect 185780 139777 185808 150350
rect 185872 140962 185900 151786
rect 185950 143440 186006 143449
rect 185950 143375 186006 143384
rect 185860 140956 185912 140962
rect 185860 140898 185912 140904
rect 185858 140584 185914 140593
rect 185964 140570 185992 143375
rect 185914 140542 185992 140570
rect 185858 140519 185914 140528
rect 185872 139890 185900 140519
rect 185872 139862 185932 139890
rect 185766 139768 185822 139777
rect 185766 139703 185822 139712
rect 184662 139496 184718 139505
rect 182822 139431 182878 139440
rect 183284 139460 183336 139466
rect 181904 139402 181956 139408
rect 184662 139431 184718 139440
rect 183284 139402 183336 139408
rect 126428 139334 126480 139340
rect 126702 139360 126758 139369
rect 126150 139295 126206 139304
rect 126702 139295 126758 139304
rect 128266 139360 128322 139369
rect 128266 139295 128322 139304
rect 132222 139360 132278 139369
rect 132222 139295 132278 139304
rect 133050 139360 133106 139369
rect 133050 139295 133106 139304
rect 145746 139360 145802 139369
rect 145746 139295 145802 139304
rect 150898 139360 150954 139369
rect 150898 139295 150954 139304
rect 154026 139360 154082 139369
rect 154026 139295 154082 139304
rect 155682 139360 155738 139369
rect 155682 139295 155738 139304
rect 155866 139360 155922 139369
rect 155866 139295 155922 139304
rect 157062 139360 157118 139369
rect 157062 139295 157118 139304
rect 159546 139360 159602 139369
rect 159546 139295 159602 139304
rect 159730 139360 159786 139369
rect 159730 139295 159786 139304
rect 178406 139360 178462 139369
rect 178406 139295 178462 139304
rect 178866 139360 178922 139369
rect 178866 139295 178922 139304
rect 180246 139360 180302 139369
rect 180246 139295 180302 139304
rect 179326 80744 179382 80753
rect 130016 80708 130068 80714
rect 130016 80650 130068 80656
rect 131672 80708 131724 80714
rect 131672 80650 131724 80656
rect 131856 80708 131908 80714
rect 179326 80679 179382 80688
rect 179602 80744 179658 80753
rect 179602 80679 179658 80688
rect 179878 80744 179934 80753
rect 179878 80679 179934 80688
rect 131856 80650 131908 80656
rect 129464 79824 129516 79830
rect 129464 79766 129516 79772
rect 124128 79620 124180 79626
rect 124128 79562 124180 79568
rect 124140 79393 124168 79562
rect 125600 79552 125652 79558
rect 125600 79494 125652 79500
rect 124126 79384 124182 79393
rect 124126 79319 124182 79328
rect 125612 77246 125640 79494
rect 126244 79484 126296 79490
rect 126244 79426 126296 79432
rect 124864 77240 124916 77246
rect 124864 77182 124916 77188
rect 125600 77240 125652 77246
rect 125600 77182 125652 77188
rect 123850 72519 123906 72528
rect 123944 72548 123996 72554
rect 123944 72490 123996 72496
rect 122104 71732 122156 71738
rect 122104 71674 122156 71680
rect 122840 71732 122892 71738
rect 122840 71674 122892 71680
rect 123300 71732 123352 71738
rect 123300 71674 123352 71680
rect 122012 70100 122064 70106
rect 122012 70042 122064 70048
rect 119804 69692 119856 69698
rect 119804 69634 119856 69640
rect 118332 69012 118384 69018
rect 118332 68954 118384 68960
rect 120080 68536 120132 68542
rect 120080 68478 120132 68484
rect 118608 68468 118660 68474
rect 118608 68410 118660 68416
rect 118620 67454 118648 68410
rect 118608 67448 118660 67454
rect 118608 67390 118660 67396
rect 118620 66858 118648 67390
rect 118620 66830 118740 66858
rect 117412 3868 117464 3874
rect 117412 3810 117464 3816
rect 118712 3398 118740 66830
rect 120092 16574 120120 68478
rect 120092 16546 120672 16574
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 118792 2916 118844 2922
rect 118792 2858 118844 2864
rect 118804 480 118832 2858
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122116 2922 122144 71674
rect 124680 3936 124732 3942
rect 124680 3878 124732 3884
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 122288 3120 122340 3126
rect 122288 3062 122340 3068
rect 122104 2916 122156 2922
rect 122104 2858 122156 2864
rect 122300 480 122328 3062
rect 123496 480 123524 3470
rect 124692 480 124720 3878
rect 124876 3126 124904 77182
rect 126256 76498 126284 79426
rect 129476 77858 129504 79766
rect 130028 78169 130056 80650
rect 130752 80368 130804 80374
rect 130752 80310 130804 80316
rect 130934 80336 130990 80345
rect 130764 80102 130792 80310
rect 130934 80271 130990 80280
rect 130752 80096 130804 80102
rect 130804 80044 130884 80054
rect 130752 80038 130884 80044
rect 130660 80028 130712 80034
rect 130764 80026 130884 80038
rect 130660 79970 130712 79976
rect 130476 79960 130528 79966
rect 130198 79928 130254 79937
rect 130476 79902 130528 79908
rect 130198 79863 130254 79872
rect 130106 79384 130162 79393
rect 130106 79319 130162 79328
rect 130120 78810 130148 79319
rect 130108 78804 130160 78810
rect 130108 78746 130160 78752
rect 130212 78198 130240 79863
rect 130488 78470 130516 79902
rect 130476 78464 130528 78470
rect 130476 78406 130528 78412
rect 130200 78192 130252 78198
rect 130014 78160 130070 78169
rect 130200 78134 130252 78140
rect 130014 78095 130070 78104
rect 129832 78056 129884 78062
rect 129832 77998 129884 78004
rect 129464 77852 129516 77858
rect 129464 77794 129516 77800
rect 129556 77852 129608 77858
rect 129556 77794 129608 77800
rect 126244 76492 126296 76498
rect 126244 76434 126296 76440
rect 126256 71806 126284 76434
rect 128912 72004 128964 72010
rect 128912 71946 128964 71952
rect 124956 71800 125008 71806
rect 124956 71742 125008 71748
rect 126244 71800 126296 71806
rect 126244 71742 126296 71748
rect 127348 71800 127400 71806
rect 127348 71742 127400 71748
rect 124968 3534 124996 71742
rect 127360 71602 127388 71742
rect 127440 71732 127492 71738
rect 127440 71674 127492 71680
rect 127452 71618 127480 71674
rect 127452 71602 127848 71618
rect 127348 71596 127400 71602
rect 127452 71596 127860 71602
rect 127452 71590 127808 71596
rect 127348 71538 127400 71544
rect 127808 71538 127860 71544
rect 128360 70916 128412 70922
rect 128360 70858 128412 70864
rect 127624 4140 127676 4146
rect 127624 4082 127676 4088
rect 125876 3868 125928 3874
rect 125876 3810 125928 3816
rect 124956 3528 125008 3534
rect 124956 3470 125008 3476
rect 124864 3120 124916 3126
rect 124864 3062 124916 3068
rect 125888 480 125916 3810
rect 127636 3738 127664 4082
rect 127624 3732 127676 3738
rect 127624 3674 127676 3680
rect 127716 3664 127768 3670
rect 127900 3664 127952 3670
rect 127768 3612 127900 3618
rect 127716 3606 127952 3612
rect 127728 3590 127940 3606
rect 128176 3596 128228 3602
rect 128176 3538 128228 3544
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 126992 480 127020 3470
rect 128188 480 128216 3538
rect 128372 490 128400 70858
rect 128924 70145 128952 71946
rect 129568 70854 129596 77794
rect 129738 75848 129794 75857
rect 129738 75783 129794 75792
rect 129556 70848 129608 70854
rect 129556 70790 129608 70796
rect 128910 70136 128966 70145
rect 128910 70071 128966 70080
rect 128452 69692 128504 69698
rect 128452 69634 128504 69640
rect 128464 3534 128492 69634
rect 128452 3528 128504 3534
rect 128452 3470 128504 3476
rect 129752 3482 129780 75783
rect 129844 3738 129872 77998
rect 130028 75138 130056 78095
rect 130200 77376 130252 77382
rect 130200 77318 130252 77324
rect 130016 75132 130068 75138
rect 130016 75074 130068 75080
rect 129924 72412 129976 72418
rect 129924 72354 129976 72360
rect 129936 3874 129964 72354
rect 130212 69630 130240 77318
rect 130292 76968 130344 76974
rect 130292 76910 130344 76916
rect 130304 76401 130332 76910
rect 130384 76900 130436 76906
rect 130384 76842 130436 76848
rect 130396 76537 130424 76842
rect 130382 76528 130438 76537
rect 130382 76463 130438 76472
rect 130290 76392 130346 76401
rect 130290 76327 130346 76336
rect 130382 75984 130438 75993
rect 130382 75919 130438 75928
rect 130200 69624 130252 69630
rect 130200 69566 130252 69572
rect 129924 3868 129976 3874
rect 129924 3810 129976 3816
rect 129832 3732 129884 3738
rect 129832 3674 129884 3680
rect 130396 3602 130424 75919
rect 130672 72758 130700 79970
rect 130856 78656 130884 80026
rect 130764 78628 130884 78656
rect 130660 72752 130712 72758
rect 130660 72694 130712 72700
rect 130764 3874 130792 78628
rect 130842 78568 130898 78577
rect 130842 78503 130844 78512
rect 130896 78503 130898 78512
rect 130844 78474 130896 78480
rect 130856 4010 130884 78474
rect 130844 4004 130896 4010
rect 130844 3946 130896 3952
rect 130752 3868 130804 3874
rect 130752 3810 130804 3816
rect 130948 3602 130976 80271
rect 131580 80164 131632 80170
rect 131580 80106 131632 80112
rect 131028 77920 131080 77926
rect 131028 77862 131080 77868
rect 131040 75857 131068 77862
rect 131212 77648 131264 77654
rect 131212 77590 131264 77596
rect 131026 75848 131082 75857
rect 131026 75783 131082 75792
rect 131028 75132 131080 75138
rect 131028 75074 131080 75080
rect 131040 68610 131068 75074
rect 131028 68604 131080 68610
rect 131028 68546 131080 68552
rect 131224 16574 131252 77590
rect 131592 70038 131620 80106
rect 131684 80102 131712 80650
rect 131868 80306 131896 80650
rect 178776 80640 178828 80646
rect 131946 80608 132002 80617
rect 131946 80543 132002 80552
rect 177762 80608 177818 80617
rect 178776 80582 178828 80588
rect 177762 80543 177818 80552
rect 131856 80300 131908 80306
rect 131856 80242 131908 80248
rect 131764 80232 131816 80238
rect 131764 80174 131816 80180
rect 131672 80096 131724 80102
rect 131672 80038 131724 80044
rect 131776 79762 131804 80174
rect 131854 80064 131910 80073
rect 131854 79999 131910 80008
rect 131764 79756 131816 79762
rect 131764 79698 131816 79704
rect 131868 79422 131896 79999
rect 131764 79416 131816 79422
rect 131764 79358 131816 79364
rect 131856 79416 131908 79422
rect 131856 79358 131908 79364
rect 131776 77586 131804 79358
rect 131856 78736 131908 78742
rect 131856 78678 131908 78684
rect 131868 78062 131896 78678
rect 131856 78056 131908 78062
rect 131856 77998 131908 78004
rect 131960 77790 131988 80543
rect 177776 80510 177804 80543
rect 177764 80504 177816 80510
rect 177764 80446 177816 80452
rect 178130 80472 178186 80481
rect 178130 80407 178186 80416
rect 178040 80368 178092 80374
rect 178040 80310 178092 80316
rect 132052 80022 132388 80050
rect 132052 78674 132080 80022
rect 132132 79892 132184 79898
rect 132132 79834 132184 79840
rect 132144 79665 132172 79834
rect 132222 79792 132278 79801
rect 132466 79744 132494 80036
rect 132558 79971 132586 80036
rect 132544 79962 132600 79971
rect 132650 79966 132678 80036
rect 132544 79897 132600 79906
rect 132638 79960 132690 79966
rect 132742 79937 132770 80036
rect 132834 79966 132862 80036
rect 132822 79960 132874 79966
rect 132638 79902 132690 79908
rect 132728 79928 132784 79937
rect 132822 79902 132874 79908
rect 132926 79898 132954 80036
rect 133018 79971 133046 80036
rect 133004 79962 133060 79971
rect 133110 79966 133138 80036
rect 132728 79863 132784 79872
rect 132914 79892 132966 79898
rect 133004 79897 133060 79906
rect 133098 79960 133150 79966
rect 133098 79902 133150 79908
rect 133202 79898 133230 80036
rect 133294 79966 133322 80036
rect 133386 79966 133414 80036
rect 133478 79966 133506 80036
rect 133570 79966 133598 80036
rect 133282 79960 133334 79966
rect 133282 79902 133334 79908
rect 133374 79960 133426 79966
rect 133374 79902 133426 79908
rect 133466 79960 133518 79966
rect 133466 79902 133518 79908
rect 133558 79960 133610 79966
rect 133558 79902 133610 79908
rect 132914 79834 132966 79840
rect 133190 79892 133242 79898
rect 133190 79834 133242 79840
rect 133512 79824 133564 79830
rect 132278 79736 132494 79744
rect 132222 79727 132494 79736
rect 132682 79792 132738 79801
rect 133326 79792 133382 79801
rect 132682 79727 132738 79736
rect 133144 79756 133196 79762
rect 132236 79716 132494 79727
rect 132130 79656 132186 79665
rect 132130 79591 132186 79600
rect 132040 78668 132092 78674
rect 132040 78610 132092 78616
rect 131948 77784 132000 77790
rect 131948 77726 132000 77732
rect 131764 77580 131816 77586
rect 131764 77522 131816 77528
rect 131776 77330 131804 77522
rect 131684 77302 131804 77330
rect 131684 75993 131712 77302
rect 131670 75984 131726 75993
rect 131670 75919 131726 75928
rect 131580 70032 131632 70038
rect 131580 69974 131632 69980
rect 132144 67634 132172 79591
rect 132236 68241 132264 79716
rect 132408 79552 132460 79558
rect 132408 79494 132460 79500
rect 132316 79348 132368 79354
rect 132316 79290 132368 79296
rect 132328 77654 132356 79290
rect 132316 77648 132368 77654
rect 132316 77590 132368 77596
rect 132420 75274 132448 79494
rect 132592 78396 132644 78402
rect 132592 78338 132644 78344
rect 132604 78169 132632 78338
rect 132590 78160 132646 78169
rect 132590 78095 132646 78104
rect 132696 78044 132724 79727
rect 133512 79766 133564 79772
rect 133326 79727 133382 79736
rect 133420 79756 133472 79762
rect 133144 79698 133196 79704
rect 133052 79620 133104 79626
rect 133052 79562 133104 79568
rect 133064 78577 133092 79562
rect 132866 78568 132922 78577
rect 132866 78503 132922 78512
rect 133050 78568 133106 78577
rect 133050 78503 133106 78512
rect 132604 78016 132724 78044
rect 132500 77988 132552 77994
rect 132500 77930 132552 77936
rect 132408 75268 132460 75274
rect 132408 75210 132460 75216
rect 132512 72418 132540 77930
rect 132500 72412 132552 72418
rect 132500 72354 132552 72360
rect 132222 68232 132278 68241
rect 132222 68167 132278 68176
rect 131776 67606 132172 67634
rect 132604 67634 132632 78016
rect 132776 77308 132828 77314
rect 132776 77250 132828 77256
rect 132684 76968 132736 76974
rect 132788 76956 132816 77250
rect 132736 76928 132816 76956
rect 132684 76910 132736 76916
rect 132776 76696 132828 76702
rect 132776 76638 132828 76644
rect 132788 76362 132816 76638
rect 132776 76356 132828 76362
rect 132776 76298 132828 76304
rect 132880 67634 132908 78503
rect 132958 78432 133014 78441
rect 132958 78367 133014 78376
rect 132972 78169 133000 78367
rect 132958 78160 133014 78169
rect 132958 78095 133014 78104
rect 133156 77330 133184 79698
rect 133340 79694 133368 79727
rect 133420 79698 133472 79704
rect 133328 79688 133380 79694
rect 133328 79630 133380 79636
rect 133236 79348 133288 79354
rect 133236 79290 133288 79296
rect 133064 77302 133184 77330
rect 132960 74792 133012 74798
rect 132960 74734 133012 74740
rect 132604 67606 132724 67634
rect 131224 16546 131344 16574
rect 130384 3596 130436 3602
rect 130384 3538 130436 3544
rect 130936 3596 130988 3602
rect 130936 3538 130988 3544
rect 129752 3454 130608 3482
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128372 462 128952 490
rect 130580 480 130608 3454
rect 128924 354 128952 462
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 131776 3398 131804 67606
rect 132696 64874 132724 67606
rect 132512 64846 132724 64874
rect 132788 67606 132908 67634
rect 132512 64190 132540 64846
rect 132500 64184 132552 64190
rect 132500 64126 132552 64132
rect 132788 63510 132816 67606
rect 132972 64874 133000 74734
rect 132880 64846 133000 64874
rect 132776 63504 132828 63510
rect 132776 63446 132828 63452
rect 132880 40730 132908 64846
rect 133064 53786 133092 77302
rect 133144 77240 133196 77246
rect 133144 77182 133196 77188
rect 133156 77042 133184 77182
rect 133144 77036 133196 77042
rect 133144 76978 133196 76984
rect 133144 76492 133196 76498
rect 133144 76434 133196 76440
rect 133156 76226 133184 76434
rect 133144 76220 133196 76226
rect 133144 76162 133196 76168
rect 133248 72010 133276 79290
rect 133328 76968 133380 76974
rect 133328 76910 133380 76916
rect 133340 76498 133368 76910
rect 133328 76492 133380 76498
rect 133328 76434 133380 76440
rect 133236 72004 133288 72010
rect 133236 71946 133288 71952
rect 133432 56574 133460 79698
rect 133524 76673 133552 79766
rect 133662 79642 133690 80036
rect 133754 79966 133782 80036
rect 133846 79966 133874 80036
rect 133938 79966 133966 80036
rect 133742 79960 133794 79966
rect 133742 79902 133794 79908
rect 133834 79960 133886 79966
rect 133926 79960 133978 79966
rect 133834 79902 133886 79908
rect 133924 79928 133926 79937
rect 133978 79928 133980 79937
rect 134030 79898 134058 80036
rect 134122 79966 134150 80036
rect 134110 79960 134162 79966
rect 134110 79902 134162 79908
rect 134214 79898 134242 80036
rect 134306 79898 134334 80036
rect 134398 79966 134426 80036
rect 134386 79960 134438 79966
rect 134386 79902 134438 79908
rect 133924 79863 133980 79872
rect 134018 79892 134070 79898
rect 134018 79834 134070 79840
rect 134202 79892 134254 79898
rect 134202 79834 134254 79840
rect 134294 79892 134346 79898
rect 134294 79834 134346 79840
rect 133742 79824 133794 79830
rect 134490 79812 134518 80036
rect 134582 79966 134610 80036
rect 134570 79960 134622 79966
rect 134570 79902 134622 79908
rect 134674 79812 134702 80036
rect 134766 79898 134794 80036
rect 134858 79937 134886 80036
rect 134950 79966 134978 80036
rect 135042 79971 135070 80036
rect 134938 79960 134990 79966
rect 134844 79928 134900 79937
rect 134754 79892 134806 79898
rect 134938 79902 134990 79908
rect 135028 79962 135084 79971
rect 135028 79897 135084 79906
rect 134844 79863 134900 79872
rect 134754 79834 134806 79840
rect 135134 79835 135162 80036
rect 135226 79966 135254 80036
rect 135318 79966 135346 80036
rect 135410 79971 135438 80036
rect 135214 79960 135266 79966
rect 135214 79902 135266 79908
rect 135306 79960 135358 79966
rect 135306 79902 135358 79908
rect 135396 79962 135452 79971
rect 135396 79897 135452 79906
rect 133794 79784 133920 79812
rect 134490 79801 134564 79812
rect 134490 79792 134578 79801
rect 134490 79784 134522 79792
rect 133742 79766 133794 79772
rect 133616 79614 133690 79642
rect 133788 79688 133840 79694
rect 133788 79630 133840 79636
rect 133616 77382 133644 79614
rect 133696 78668 133748 78674
rect 133696 78610 133748 78616
rect 133604 77376 133656 77382
rect 133604 77318 133656 77324
rect 133604 76900 133656 76906
rect 133604 76842 133656 76848
rect 133510 76664 133566 76673
rect 133510 76599 133566 76608
rect 133524 74798 133552 76599
rect 133616 76537 133644 76842
rect 133602 76528 133658 76537
rect 133602 76463 133658 76472
rect 133512 74792 133564 74798
rect 133512 74734 133564 74740
rect 133708 67634 133736 78610
rect 133800 74186 133828 79630
rect 133892 78674 133920 79784
rect 134248 79756 134300 79762
rect 134522 79727 134578 79736
rect 134628 79784 134702 79812
rect 135120 79826 135176 79835
rect 134248 79698 134300 79704
rect 134156 79688 134208 79694
rect 134156 79630 134208 79636
rect 134064 79620 134116 79626
rect 134064 79562 134116 79568
rect 133880 78668 133932 78674
rect 133880 78610 133932 78616
rect 134076 78606 134104 79562
rect 134064 78600 134116 78606
rect 134064 78542 134116 78548
rect 133880 78532 133932 78538
rect 133880 78474 133932 78480
rect 133892 78198 133920 78474
rect 133880 78192 133932 78198
rect 133880 78134 133932 78140
rect 134062 77480 134118 77489
rect 134062 77415 134064 77424
rect 134116 77415 134118 77424
rect 134064 77386 134116 77392
rect 134064 76832 134116 76838
rect 134064 76774 134116 76780
rect 134076 76401 134104 76774
rect 134062 76392 134118 76401
rect 134062 76327 134118 76336
rect 134168 74225 134196 79630
rect 134260 77058 134288 79698
rect 134432 79688 134484 79694
rect 134432 79630 134484 79636
rect 134340 79620 134392 79626
rect 134340 79562 134392 79568
rect 134352 77194 134380 79562
rect 134444 77858 134472 79630
rect 134524 79552 134576 79558
rect 134524 79494 134576 79500
rect 134432 77852 134484 77858
rect 134432 77794 134484 77800
rect 134536 77217 134564 79494
rect 134522 77208 134578 77217
rect 134352 77166 134472 77194
rect 134260 77030 134380 77058
rect 134246 76664 134302 76673
rect 134246 76599 134302 76608
rect 134154 74216 134210 74225
rect 133788 74180 133840 74186
rect 134154 74151 134210 74160
rect 133788 74122 133840 74128
rect 134156 73976 134208 73982
rect 134156 73918 134208 73924
rect 133616 67606 133736 67634
rect 133616 60722 133644 67606
rect 133604 60716 133656 60722
rect 133604 60658 133656 60664
rect 133420 56568 133472 56574
rect 133420 56510 133472 56516
rect 133052 53780 133104 53786
rect 133052 53722 133104 53728
rect 132868 40724 132920 40730
rect 132868 40666 132920 40672
rect 134168 7614 134196 73918
rect 134260 39370 134288 76599
rect 134352 72282 134380 77030
rect 134340 72276 134392 72282
rect 134340 72218 134392 72224
rect 134340 72140 134392 72146
rect 134340 72082 134392 72088
rect 134352 66230 134380 72082
rect 134444 71670 134472 77166
rect 134522 77143 134578 77152
rect 134524 76696 134576 76702
rect 134524 76638 134576 76644
rect 134432 71664 134484 71670
rect 134432 71606 134484 71612
rect 134340 66224 134392 66230
rect 134340 66166 134392 66172
rect 134248 39364 134300 39370
rect 134248 39306 134300 39312
rect 134156 7608 134208 7614
rect 134156 7550 134208 7556
rect 134536 4146 134564 76638
rect 134628 73982 134656 79784
rect 135352 79824 135404 79830
rect 135120 79761 135176 79770
rect 135258 79792 135314 79801
rect 135502 79812 135530 80036
rect 135352 79766 135404 79772
rect 135456 79784 135530 79812
rect 135258 79727 135314 79736
rect 135168 79688 135220 79694
rect 135074 79656 135130 79665
rect 134708 79620 134760 79626
rect 135168 79630 135220 79636
rect 135074 79591 135130 79600
rect 134708 79562 134760 79568
rect 134720 75993 134748 79562
rect 135088 79558 135116 79591
rect 135076 79552 135128 79558
rect 135076 79494 135128 79500
rect 134706 75984 134762 75993
rect 134706 75919 134762 75928
rect 134616 73976 134668 73982
rect 134616 73918 134668 73924
rect 135180 72146 135208 79630
rect 135272 76566 135300 79727
rect 135260 76560 135312 76566
rect 135260 76502 135312 76508
rect 135364 75857 135392 79766
rect 135456 75993 135484 79784
rect 135594 79744 135622 80036
rect 135686 79830 135714 80036
rect 135778 79830 135806 80036
rect 135674 79824 135726 79830
rect 135674 79766 135726 79772
rect 135766 79824 135818 79830
rect 135766 79766 135818 79772
rect 135548 79716 135622 79744
rect 135870 79744 135898 80036
rect 135962 79898 135990 80036
rect 135950 79892 136002 79898
rect 135950 79834 136002 79840
rect 136054 79778 136082 80036
rect 136146 79966 136174 80036
rect 136134 79960 136186 79966
rect 136134 79902 136186 79908
rect 136238 79898 136266 80036
rect 136330 79966 136358 80036
rect 136422 79971 136450 80036
rect 136318 79960 136370 79966
rect 136318 79902 136370 79908
rect 136408 79962 136464 79971
rect 136226 79892 136278 79898
rect 136408 79897 136464 79906
rect 136226 79834 136278 79840
rect 136364 79824 136416 79830
rect 136054 79750 136128 79778
rect 136514 79812 136542 80036
rect 136416 79784 136542 79812
rect 136364 79766 136416 79772
rect 135870 79716 135944 79744
rect 135548 79354 135576 79716
rect 135720 79688 135772 79694
rect 135718 79656 135720 79665
rect 135772 79656 135774 79665
rect 135628 79620 135680 79626
rect 135718 79591 135774 79600
rect 135628 79562 135680 79568
rect 135536 79348 135588 79354
rect 135536 79290 135588 79296
rect 135640 78656 135668 79562
rect 135548 78628 135668 78656
rect 135442 75984 135498 75993
rect 135442 75919 135498 75928
rect 135350 75848 135406 75857
rect 135350 75783 135406 75792
rect 135444 75608 135496 75614
rect 135444 75550 135496 75556
rect 135456 74934 135484 75550
rect 135444 74928 135496 74934
rect 135444 74870 135496 74876
rect 135168 72140 135220 72146
rect 135168 72082 135220 72088
rect 135260 68604 135312 68610
rect 135260 68546 135312 68552
rect 134524 4140 134576 4146
rect 134524 4082 134576 4088
rect 131764 3392 131816 3398
rect 131764 3334 131816 3340
rect 134156 3120 134208 3126
rect 134156 3062 134208 3068
rect 132960 3052 133012 3058
rect 132960 2994 133012 3000
rect 132972 480 133000 2994
rect 134168 480 134196 3062
rect 135272 480 135300 68546
rect 135352 61940 135404 61946
rect 135352 61882 135404 61888
rect 135364 16574 135392 61882
rect 135456 35222 135484 74870
rect 135548 74118 135576 78628
rect 135626 78568 135682 78577
rect 135626 78503 135682 78512
rect 135536 74112 135588 74118
rect 135536 74054 135588 74060
rect 135444 35216 135496 35222
rect 135444 35158 135496 35164
rect 135548 31074 135576 74054
rect 135640 37942 135668 78503
rect 135732 61402 135760 79591
rect 135812 79552 135864 79558
rect 135812 79494 135864 79500
rect 135824 77897 135852 79494
rect 135810 77888 135866 77897
rect 135810 77823 135866 77832
rect 135824 76634 135852 77823
rect 135812 76628 135864 76634
rect 135812 76570 135864 76576
rect 135916 75993 135944 79716
rect 135996 79688 136048 79694
rect 135996 79630 136048 79636
rect 136008 78305 136036 79630
rect 135994 78296 136050 78305
rect 135994 78231 136050 78240
rect 135902 75984 135958 75993
rect 135902 75919 135958 75928
rect 135812 75268 135864 75274
rect 135812 75210 135864 75216
rect 135824 62082 135852 75210
rect 136008 71058 136036 78231
rect 136100 77518 136128 79750
rect 136272 79756 136324 79762
rect 136606 79744 136634 80036
rect 136698 79966 136726 80036
rect 136790 79971 136818 80036
rect 136686 79960 136738 79966
rect 136686 79902 136738 79908
rect 136776 79962 136832 79971
rect 136776 79897 136832 79906
rect 136272 79698 136324 79704
rect 136560 79716 136634 79744
rect 136732 79756 136784 79762
rect 136180 79688 136232 79694
rect 136180 79630 136232 79636
rect 136088 77512 136140 77518
rect 136088 77454 136140 77460
rect 136192 75256 136220 79630
rect 136100 75228 136220 75256
rect 135996 71052 136048 71058
rect 135996 70994 136048 71000
rect 136100 68814 136128 75228
rect 136284 70394 136312 79698
rect 136362 79656 136418 79665
rect 136362 79591 136418 79600
rect 136376 75274 136404 79591
rect 136456 79552 136508 79558
rect 136456 79494 136508 79500
rect 136364 75268 136416 75274
rect 136364 75210 136416 75216
rect 136468 73710 136496 79494
rect 136560 74934 136588 79716
rect 136882 79744 136910 80036
rect 136974 79812 137002 80036
rect 137066 79971 137094 80036
rect 137052 79962 137108 79971
rect 137158 79966 137186 80036
rect 137052 79897 137108 79906
rect 137146 79960 137198 79966
rect 137146 79902 137198 79908
rect 136974 79784 137048 79812
rect 136732 79698 136784 79704
rect 136836 79716 136910 79744
rect 136548 74928 136600 74934
rect 136744 74905 136772 79698
rect 136836 77722 136864 79716
rect 136916 79620 136968 79626
rect 136916 79562 136968 79568
rect 136928 77761 136956 79562
rect 136914 77752 136970 77761
rect 136824 77716 136876 77722
rect 136914 77687 136970 77696
rect 136824 77658 136876 77664
rect 137020 77602 137048 79784
rect 137098 79792 137154 79801
rect 137250 79778 137278 80036
rect 137342 79937 137370 80036
rect 137434 79966 137462 80036
rect 137422 79960 137474 79966
rect 137328 79928 137384 79937
rect 137422 79902 137474 79908
rect 137328 79863 137384 79872
rect 137098 79727 137100 79736
rect 137152 79727 137154 79736
rect 137204 79750 137278 79778
rect 137342 79778 137370 79863
rect 137526 79812 137554 80036
rect 137480 79784 137554 79812
rect 137342 79750 137416 79778
rect 137100 79698 137152 79704
rect 137100 78464 137152 78470
rect 137100 78406 137152 78412
rect 137112 77994 137140 78406
rect 137100 77988 137152 77994
rect 137100 77930 137152 77936
rect 137100 77716 137152 77722
rect 137100 77658 137152 77664
rect 136928 77574 137048 77602
rect 136928 76838 136956 77574
rect 137008 77512 137060 77518
rect 137008 77454 137060 77460
rect 136916 76832 136968 76838
rect 136916 76774 136968 76780
rect 136548 74870 136600 74876
rect 136730 74896 136786 74905
rect 136730 74831 136786 74840
rect 136456 73704 136508 73710
rect 136456 73646 136508 73652
rect 136824 70984 136876 70990
rect 136824 70926 136876 70932
rect 136192 70366 136312 70394
rect 136088 68808 136140 68814
rect 136088 68750 136140 68756
rect 136192 67634 136220 70366
rect 136008 67606 136220 67634
rect 135812 62076 135864 62082
rect 135812 62018 135864 62024
rect 135720 61396 135772 61402
rect 135720 61338 135772 61344
rect 136008 59362 136036 67606
rect 135996 59356 136048 59362
rect 135996 59298 136048 59304
rect 135628 37936 135680 37942
rect 135628 37878 135680 37884
rect 135536 31068 135588 31074
rect 135536 31010 135588 31016
rect 135364 16546 136496 16574
rect 136468 480 136496 16546
rect 136836 3126 136864 70926
rect 137020 55962 137048 77454
rect 137112 70922 137140 77658
rect 137100 70916 137152 70922
rect 137100 70858 137152 70864
rect 137204 64870 137232 79750
rect 137284 79688 137336 79694
rect 137284 79630 137336 79636
rect 137296 78305 137324 79630
rect 137282 78296 137338 78305
rect 137282 78231 137338 78240
rect 137192 64864 137244 64870
rect 137192 64806 137244 64812
rect 137008 55956 137060 55962
rect 137008 55898 137060 55904
rect 137296 3466 137324 78231
rect 137388 77518 137416 79750
rect 137376 77512 137428 77518
rect 137376 77454 137428 77460
rect 137480 77246 137508 79784
rect 137618 79778 137646 80036
rect 137710 79898 137738 80036
rect 137698 79892 137750 79898
rect 137698 79834 137750 79840
rect 137802 79778 137830 80036
rect 137894 79937 137922 80036
rect 137986 79966 138014 80036
rect 138078 79966 138106 80036
rect 138170 79966 138198 80036
rect 138262 79966 138290 80036
rect 138354 79971 138382 80036
rect 137974 79960 138026 79966
rect 137880 79928 137936 79937
rect 137974 79902 138026 79908
rect 138066 79960 138118 79966
rect 138066 79902 138118 79908
rect 138158 79960 138210 79966
rect 138158 79902 138210 79908
rect 138250 79960 138302 79966
rect 138250 79902 138302 79908
rect 138340 79962 138396 79971
rect 138340 79897 138396 79906
rect 137880 79863 137936 79872
rect 137894 79830 137922 79863
rect 137618 79750 137692 79778
rect 137560 79688 137612 79694
rect 137664 79665 137692 79750
rect 137756 79750 137830 79778
rect 137882 79824 137934 79830
rect 137882 79766 137934 79772
rect 138020 79824 138072 79830
rect 138020 79766 138072 79772
rect 138112 79824 138164 79830
rect 138446 79812 138474 80036
rect 138308 79801 138474 79812
rect 138112 79766 138164 79772
rect 138294 79792 138474 79801
rect 137560 79630 137612 79636
rect 137650 79656 137706 79665
rect 137572 78742 137600 79630
rect 137650 79591 137706 79600
rect 137560 78736 137612 78742
rect 137560 78678 137612 78684
rect 137560 78600 137612 78606
rect 137560 78542 137612 78548
rect 137572 78198 137600 78542
rect 137560 78192 137612 78198
rect 137560 78134 137612 78140
rect 137560 77444 137612 77450
rect 137560 77386 137612 77392
rect 137572 77353 137600 77386
rect 137558 77344 137614 77353
rect 137558 77279 137614 77288
rect 137468 77240 137520 77246
rect 137468 77182 137520 77188
rect 137664 75342 137692 79591
rect 137652 75336 137704 75342
rect 137652 75278 137704 75284
rect 137756 70394 137784 79750
rect 137836 79688 137888 79694
rect 137836 79630 137888 79636
rect 137848 72622 137876 79630
rect 137926 78568 137982 78577
rect 137926 78503 137982 78512
rect 137836 72616 137888 72622
rect 137836 72558 137888 72564
rect 137480 70366 137784 70394
rect 137480 60654 137508 70366
rect 137468 60648 137520 60654
rect 137468 60590 137520 60596
rect 137940 44878 137968 78503
rect 138032 77761 138060 79766
rect 138124 78577 138152 79766
rect 138204 79756 138256 79762
rect 138350 79784 138474 79792
rect 138538 79744 138566 80036
rect 138630 79966 138658 80036
rect 138618 79960 138670 79966
rect 138722 79937 138750 80036
rect 138618 79902 138670 79908
rect 138708 79928 138764 79937
rect 138814 79898 138842 80036
rect 138708 79863 138764 79872
rect 138802 79892 138854 79898
rect 138722 79812 138750 79863
rect 138802 79834 138854 79840
rect 138294 79727 138350 79736
rect 138204 79698 138256 79704
rect 138110 78568 138166 78577
rect 138110 78503 138166 78512
rect 138216 77976 138244 79698
rect 138308 79354 138336 79727
rect 138492 79716 138566 79744
rect 138676 79784 138750 79812
rect 138296 79348 138348 79354
rect 138296 79290 138348 79296
rect 138492 78962 138520 79716
rect 138572 79552 138624 79558
rect 138572 79494 138624 79500
rect 138400 78934 138520 78962
rect 138294 78704 138350 78713
rect 138400 78674 138428 78934
rect 138584 78792 138612 79494
rect 138492 78764 138612 78792
rect 138294 78639 138350 78648
rect 138388 78668 138440 78674
rect 138308 78266 138336 78639
rect 138388 78610 138440 78616
rect 138296 78260 138348 78266
rect 138296 78202 138348 78208
rect 138124 77948 138244 77976
rect 138018 77752 138074 77761
rect 138018 77687 138074 77696
rect 138124 77568 138152 77948
rect 138202 77888 138258 77897
rect 138202 77823 138258 77832
rect 138032 77540 138152 77568
rect 138032 75818 138060 77540
rect 138110 77480 138166 77489
rect 138110 77415 138112 77424
rect 138164 77415 138166 77424
rect 138112 77386 138164 77392
rect 138216 77353 138244 77823
rect 138294 77480 138350 77489
rect 138294 77415 138350 77424
rect 138202 77344 138258 77353
rect 138202 77279 138258 77288
rect 138020 75812 138072 75818
rect 138020 75754 138072 75760
rect 138204 71188 138256 71194
rect 138204 71130 138256 71136
rect 138112 69760 138164 69766
rect 138112 69702 138164 69708
rect 137928 44872 137980 44878
rect 137928 44814 137980 44820
rect 138020 42628 138072 42634
rect 138020 42570 138072 42576
rect 138032 6914 138060 42570
rect 138124 10334 138152 69702
rect 138112 10328 138164 10334
rect 138112 10270 138164 10276
rect 138032 6886 138152 6914
rect 137652 3664 137704 3670
rect 137652 3606 137704 3612
rect 137284 3460 137336 3466
rect 137284 3402 137336 3408
rect 136824 3120 136876 3126
rect 136824 3062 136876 3068
rect 137664 480 137692 3606
rect 138124 3482 138152 6886
rect 138216 3738 138244 71130
rect 138308 70394 138336 77415
rect 138308 70366 138428 70394
rect 138400 62898 138428 70366
rect 138492 67590 138520 78764
rect 138572 78668 138624 78674
rect 138572 78610 138624 78616
rect 138584 72894 138612 78610
rect 138676 75410 138704 79784
rect 138906 79778 138934 80036
rect 138860 79750 138934 79778
rect 138998 79778 139026 80036
rect 139090 79898 139118 80036
rect 139078 79892 139130 79898
rect 139078 79834 139130 79840
rect 139182 79778 139210 80036
rect 139274 79966 139302 80036
rect 139366 79971 139394 80036
rect 139262 79960 139314 79966
rect 139262 79902 139314 79908
rect 139352 79962 139408 79971
rect 139352 79897 139408 79906
rect 138998 79750 139072 79778
rect 138860 79540 138888 79750
rect 139044 79665 139072 79750
rect 139136 79750 139210 79778
rect 139030 79656 139086 79665
rect 139030 79591 139086 79600
rect 138768 79512 138888 79540
rect 138768 77625 138796 79512
rect 138940 79348 138992 79354
rect 138940 79290 138992 79296
rect 138848 78668 138900 78674
rect 138848 78610 138900 78616
rect 138754 77616 138810 77625
rect 138754 77551 138810 77560
rect 138664 75404 138716 75410
rect 138664 75346 138716 75352
rect 138572 72888 138624 72894
rect 138572 72830 138624 72836
rect 138860 70394 138888 78610
rect 138584 70366 138888 70394
rect 138584 69766 138612 70366
rect 138572 69760 138624 69766
rect 138572 69702 138624 69708
rect 138480 67584 138532 67590
rect 138480 67526 138532 67532
rect 138952 64874 138980 79290
rect 139044 76702 139072 79591
rect 139136 78674 139164 79750
rect 139458 79744 139486 80036
rect 139550 79937 139578 80036
rect 139642 79966 139670 80036
rect 139630 79960 139682 79966
rect 139536 79928 139592 79937
rect 139630 79902 139682 79908
rect 139536 79863 139592 79872
rect 139734 79812 139762 80036
rect 139826 79937 139854 80036
rect 139812 79928 139868 79937
rect 139812 79863 139868 79872
rect 139688 79784 139762 79812
rect 139458 79716 139532 79744
rect 139216 79688 139268 79694
rect 139214 79656 139216 79665
rect 139268 79656 139270 79665
rect 139214 79591 139270 79600
rect 139308 79620 139360 79626
rect 139308 79562 139360 79568
rect 139400 79620 139452 79626
rect 139400 79562 139452 79568
rect 139216 79552 139268 79558
rect 139216 79494 139268 79500
rect 139124 78668 139176 78674
rect 139124 78610 139176 78616
rect 139124 78396 139176 78402
rect 139124 78338 139176 78344
rect 139032 76696 139084 76702
rect 139032 76638 139084 76644
rect 139136 72962 139164 78338
rect 139124 72956 139176 72962
rect 139124 72898 139176 72904
rect 139228 71194 139256 79494
rect 139320 78402 139348 79562
rect 139308 78396 139360 78402
rect 139308 78338 139360 78344
rect 139306 78160 139362 78169
rect 139306 78095 139362 78104
rect 139320 77625 139348 78095
rect 139306 77616 139362 77625
rect 139306 77551 139362 77560
rect 139412 75886 139440 79562
rect 139400 75880 139452 75886
rect 139400 75822 139452 75828
rect 139504 75274 139532 79716
rect 139688 79665 139716 79784
rect 139918 79744 139946 80036
rect 139780 79716 139946 79744
rect 139674 79656 139730 79665
rect 139674 79591 139730 79600
rect 139780 79064 139808 79716
rect 140010 79676 140038 80036
rect 140102 79903 140130 80036
rect 140088 79894 140144 79903
rect 140088 79829 140144 79838
rect 140194 79778 140222 80036
rect 139964 79648 140038 79676
rect 140148 79750 140222 79778
rect 139860 79620 139912 79626
rect 139860 79562 139912 79568
rect 139688 79036 139808 79064
rect 139582 78976 139638 78985
rect 139582 78911 139638 78920
rect 139596 78588 139624 78911
rect 139688 78713 139716 79036
rect 139674 78704 139730 78713
rect 139674 78639 139730 78648
rect 139596 78560 139716 78588
rect 139582 77344 139638 77353
rect 139582 77279 139638 77288
rect 139492 75268 139544 75274
rect 139492 75210 139544 75216
rect 139216 71188 139268 71194
rect 139216 71130 139268 71136
rect 139492 69896 139544 69902
rect 139492 69838 139544 69844
rect 139504 69766 139532 69838
rect 139492 69760 139544 69766
rect 139492 69702 139544 69708
rect 139400 64932 139452 64938
rect 139400 64874 139452 64880
rect 138860 64846 138980 64874
rect 138388 62892 138440 62898
rect 138388 62834 138440 62840
rect 138664 55276 138716 55282
rect 138664 55218 138716 55224
rect 138204 3732 138256 3738
rect 138204 3674 138256 3680
rect 138676 3670 138704 55218
rect 138860 42090 138888 64846
rect 138848 42084 138900 42090
rect 138848 42026 138900 42032
rect 138664 3664 138716 3670
rect 138664 3606 138716 3612
rect 138124 3454 138888 3482
rect 138860 480 138888 3454
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 139412 354 139440 64874
rect 139504 3806 139532 69702
rect 139596 67046 139624 77279
rect 139584 67040 139636 67046
rect 139584 66982 139636 66988
rect 139688 66978 139716 78560
rect 139766 77752 139822 77761
rect 139766 77687 139822 77696
rect 139676 66972 139728 66978
rect 139676 66914 139728 66920
rect 139780 66910 139808 77687
rect 139872 77654 139900 79562
rect 139860 77648 139912 77654
rect 139860 77590 139912 77596
rect 139964 75682 139992 79648
rect 140044 79552 140096 79558
rect 140044 79494 140096 79500
rect 140056 78810 140084 79494
rect 140044 78804 140096 78810
rect 140044 78746 140096 78752
rect 140148 76294 140176 79750
rect 140286 79744 140314 80036
rect 140378 79966 140406 80036
rect 140470 79966 140498 80036
rect 140562 79966 140590 80036
rect 140366 79960 140418 79966
rect 140366 79902 140418 79908
rect 140458 79960 140510 79966
rect 140458 79902 140510 79908
rect 140550 79960 140602 79966
rect 140654 79937 140682 80036
rect 140550 79902 140602 79908
rect 140640 79928 140696 79937
rect 140640 79863 140696 79872
rect 140412 79824 140464 79830
rect 140746 79812 140774 80036
rect 140838 79937 140866 80036
rect 140824 79928 140880 79937
rect 140824 79863 140880 79872
rect 140412 79766 140464 79772
rect 140608 79784 140774 79812
rect 140286 79716 140360 79744
rect 140228 79620 140280 79626
rect 140228 79562 140280 79568
rect 140136 76288 140188 76294
rect 140136 76230 140188 76236
rect 139952 75676 140004 75682
rect 139952 75618 140004 75624
rect 140240 70394 140268 79562
rect 140332 76378 140360 79716
rect 140424 76498 140452 79766
rect 140504 78940 140556 78946
rect 140504 78882 140556 78888
rect 140516 78674 140544 78882
rect 140504 78668 140556 78674
rect 140504 78610 140556 78616
rect 140412 76492 140464 76498
rect 140412 76434 140464 76440
rect 140332 76350 140452 76378
rect 140320 75268 140372 75274
rect 140320 75210 140372 75216
rect 139872 70366 140268 70394
rect 139872 67522 139900 70366
rect 140332 69766 140360 75210
rect 140424 71126 140452 76350
rect 140608 71466 140636 79784
rect 140930 79744 140958 80036
rect 141022 79898 141050 80036
rect 141010 79892 141062 79898
rect 141010 79834 141062 79840
rect 141114 79744 141142 80036
rect 141206 79801 141234 80036
rect 140930 79716 141004 79744
rect 140778 79656 140834 79665
rect 140778 79591 140834 79600
rect 140688 79552 140740 79558
rect 140688 79494 140740 79500
rect 140700 78985 140728 79494
rect 140686 78976 140742 78985
rect 140686 78911 140742 78920
rect 140596 71460 140648 71466
rect 140596 71402 140648 71408
rect 140412 71120 140464 71126
rect 140412 71062 140464 71068
rect 140320 69760 140372 69766
rect 140320 69702 140372 69708
rect 140792 68338 140820 79591
rect 140872 79552 140924 79558
rect 140872 79494 140924 79500
rect 140884 78985 140912 79494
rect 140870 78976 140926 78985
rect 140870 78911 140926 78920
rect 140976 78742 141004 79716
rect 141068 79716 141142 79744
rect 141192 79792 141248 79801
rect 141192 79727 141248 79736
rect 140964 78736 141016 78742
rect 140964 78678 141016 78684
rect 140964 78396 141016 78402
rect 140964 78338 141016 78344
rect 140870 77480 140926 77489
rect 140870 77415 140926 77424
rect 140780 68332 140832 68338
rect 140780 68274 140832 68280
rect 139860 67516 139912 67522
rect 139860 67458 139912 67464
rect 139768 66904 139820 66910
rect 139768 66846 139820 66852
rect 139872 8974 139900 67458
rect 140780 66292 140832 66298
rect 140780 66234 140832 66240
rect 139860 8968 139912 8974
rect 139860 8910 139912 8916
rect 139492 3800 139544 3806
rect 139492 3742 139544 3748
rect 140792 1306 140820 66234
rect 140884 3942 140912 77415
rect 140976 68406 141004 78338
rect 141068 76362 141096 79716
rect 141298 79676 141326 80036
rect 141390 79812 141418 80036
rect 141482 79966 141510 80036
rect 141574 79966 141602 80036
rect 141470 79960 141522 79966
rect 141470 79902 141522 79908
rect 141562 79960 141614 79966
rect 141562 79902 141614 79908
rect 141666 79898 141694 80036
rect 141758 79937 141786 80036
rect 141744 79928 141800 79937
rect 141654 79892 141706 79898
rect 141850 79898 141878 80036
rect 141744 79863 141800 79872
rect 141838 79892 141890 79898
rect 141654 79834 141706 79840
rect 141390 79784 141602 79812
rect 141574 79778 141602 79784
rect 141574 79750 141648 79778
rect 141160 79648 141326 79676
rect 141422 79656 141478 79665
rect 141056 76356 141108 76362
rect 141056 76298 141108 76304
rect 141160 72690 141188 79648
rect 141422 79591 141424 79600
rect 141476 79591 141478 79600
rect 141424 79562 141476 79568
rect 141240 79552 141292 79558
rect 141240 79494 141292 79500
rect 141148 72684 141200 72690
rect 141148 72626 141200 72632
rect 141252 68474 141280 79494
rect 141332 79212 141384 79218
rect 141332 79154 141384 79160
rect 141344 78946 141372 79154
rect 141332 78940 141384 78946
rect 141332 78882 141384 78888
rect 141332 78736 141384 78742
rect 141332 78678 141384 78684
rect 141344 77217 141372 78678
rect 141436 78402 141464 79562
rect 141424 78396 141476 78402
rect 141424 78338 141476 78344
rect 141330 77208 141386 77217
rect 141330 77143 141386 77152
rect 141516 74316 141568 74322
rect 141516 74258 141568 74264
rect 141528 74186 141556 74258
rect 141516 74180 141568 74186
rect 141516 74122 141568 74128
rect 141620 72486 141648 79750
rect 141758 79744 141786 79863
rect 141838 79834 141890 79840
rect 141942 79801 141970 80036
rect 142034 79898 142062 80036
rect 142022 79892 142074 79898
rect 142022 79834 142074 79840
rect 141928 79792 141984 79801
rect 141758 79716 141832 79744
rect 142126 79744 142154 80036
rect 142218 79801 142246 80036
rect 142310 79966 142338 80036
rect 142298 79960 142350 79966
rect 142298 79902 142350 79908
rect 142402 79812 142430 80036
rect 142494 79971 142522 80036
rect 142480 79962 142536 79971
rect 142586 79966 142614 80036
rect 142480 79897 142536 79906
rect 142574 79960 142626 79966
rect 142574 79902 142626 79908
rect 141928 79727 141984 79736
rect 141698 79656 141754 79665
rect 141698 79591 141754 79600
rect 141712 76226 141740 79591
rect 141700 76220 141752 76226
rect 141700 76162 141752 76168
rect 141608 72480 141660 72486
rect 141608 72422 141660 72428
rect 141424 71664 141476 71670
rect 141424 71606 141476 71612
rect 141240 68468 141292 68474
rect 141240 68410 141292 68416
rect 140964 68400 141016 68406
rect 140964 68342 141016 68348
rect 140872 3936 140924 3942
rect 140872 3878 140924 3884
rect 141436 3058 141464 71606
rect 141804 68542 141832 79716
rect 142080 79716 142154 79744
rect 142204 79792 142260 79801
rect 142204 79727 142260 79736
rect 142356 79784 142430 79812
rect 142526 79792 142582 79801
rect 141884 79688 141936 79694
rect 141884 79630 141936 79636
rect 141976 79688 142028 79694
rect 141976 79630 142028 79636
rect 141896 77042 141924 79630
rect 141988 77489 142016 79630
rect 142080 78690 142108 79716
rect 142252 79688 142304 79694
rect 142252 79630 142304 79636
rect 142160 79484 142212 79490
rect 142160 79426 142212 79432
rect 142172 79014 142200 79426
rect 142160 79008 142212 79014
rect 142160 78950 142212 78956
rect 142080 78662 142200 78690
rect 142068 78464 142120 78470
rect 142172 78418 142200 78662
rect 142120 78412 142200 78418
rect 142068 78406 142200 78412
rect 142080 78390 142200 78406
rect 142264 77586 142292 79630
rect 142356 77722 142384 79784
rect 142678 79778 142706 80036
rect 142770 79966 142798 80036
rect 142758 79960 142810 79966
rect 142758 79902 142810 79908
rect 142862 79903 142890 80036
rect 142848 79894 142904 79903
rect 142848 79829 142904 79838
rect 142632 79762 142706 79778
rect 142526 79727 142582 79736
rect 142620 79756 142706 79762
rect 142434 79656 142490 79665
rect 142434 79591 142490 79600
rect 142344 77716 142396 77722
rect 142344 77658 142396 77664
rect 142252 77580 142304 77586
rect 142252 77522 142304 77528
rect 141974 77480 142030 77489
rect 141974 77415 142030 77424
rect 141884 77036 141936 77042
rect 141884 76978 141936 76984
rect 142252 74520 142304 74526
rect 142252 74462 142304 74468
rect 142264 73914 142292 74462
rect 142252 73908 142304 73914
rect 142252 73850 142304 73856
rect 142066 70408 142122 70417
rect 142066 70343 142122 70352
rect 141792 68536 141844 68542
rect 141792 68478 141844 68484
rect 142080 64977 142108 70343
rect 142160 69828 142212 69834
rect 142160 69770 142212 69776
rect 142172 66298 142200 69770
rect 142160 66292 142212 66298
rect 142160 66234 142212 66240
rect 142264 66178 142292 73850
rect 142448 69698 142476 79591
rect 142540 77926 142568 79727
rect 142672 79750 142706 79756
rect 142804 79756 142856 79762
rect 142620 79698 142672 79704
rect 142954 79744 142982 80036
rect 143046 79898 143074 80036
rect 143034 79892 143086 79898
rect 143034 79834 143086 79840
rect 143138 79744 143166 80036
rect 142804 79698 142856 79704
rect 142908 79716 142982 79744
rect 143092 79716 143166 79744
rect 142618 79656 142674 79665
rect 142618 79591 142674 79600
rect 142712 79620 142764 79626
rect 142632 78538 142660 79591
rect 142712 79562 142764 79568
rect 142620 78532 142672 78538
rect 142620 78474 142672 78480
rect 142620 78396 142672 78402
rect 142620 78338 142672 78344
rect 142528 77920 142580 77926
rect 142528 77862 142580 77868
rect 142632 77330 142660 78338
rect 142540 77302 142660 77330
rect 142540 73846 142568 77302
rect 142618 77208 142674 77217
rect 142618 77143 142674 77152
rect 142528 73840 142580 73846
rect 142528 73782 142580 73788
rect 142540 70718 142568 73782
rect 142528 70712 142580 70718
rect 142528 70654 142580 70660
rect 142528 69964 142580 69970
rect 142528 69906 142580 69912
rect 142436 69692 142488 69698
rect 142436 69634 142488 69640
rect 142344 68876 142396 68882
rect 142344 68818 142396 68824
rect 142172 66150 142292 66178
rect 142066 64968 142122 64977
rect 142172 64938 142200 66150
rect 142356 64954 142384 68818
rect 142066 64903 142122 64912
rect 142160 64932 142212 64938
rect 142160 64874 142212 64880
rect 142264 64926 142384 64954
rect 142066 64832 142122 64841
rect 142066 64767 142122 64776
rect 142080 55321 142108 64767
rect 142066 55312 142122 55321
rect 142066 55247 142122 55256
rect 142066 55176 142122 55185
rect 142066 55111 142122 55120
rect 142080 45665 142108 55111
rect 142066 45656 142122 45665
rect 142066 45591 142122 45600
rect 142066 45520 142122 45529
rect 142066 45455 142122 45464
rect 142080 36009 142108 45455
rect 142264 42634 142292 64926
rect 142540 64874 142568 69906
rect 142632 69834 142660 77143
rect 142620 69828 142672 69834
rect 142620 69770 142672 69776
rect 142724 68882 142752 79562
rect 142816 78962 142844 79698
rect 142908 79098 142936 79716
rect 143092 79626 143120 79716
rect 143230 79676 143258 80036
rect 143322 79937 143350 80036
rect 143414 79966 143442 80036
rect 143402 79960 143454 79966
rect 143308 79928 143364 79937
rect 143506 79937 143534 80036
rect 143402 79902 143454 79908
rect 143492 79928 143548 79937
rect 143308 79863 143364 79872
rect 143492 79863 143548 79872
rect 143598 79778 143626 80036
rect 143690 79966 143718 80036
rect 143678 79960 143730 79966
rect 143782 79937 143810 80036
rect 143678 79902 143730 79908
rect 143768 79928 143824 79937
rect 143552 79762 143626 79778
rect 143448 79756 143500 79762
rect 143448 79698 143500 79704
rect 143540 79756 143626 79762
rect 143592 79750 143626 79756
rect 143540 79698 143592 79704
rect 143184 79648 143258 79676
rect 143356 79688 143408 79694
rect 143080 79620 143132 79626
rect 143080 79562 143132 79568
rect 143080 79484 143132 79490
rect 143080 79426 143132 79432
rect 142988 79416 143040 79422
rect 142988 79358 143040 79364
rect 143000 79218 143028 79358
rect 142988 79212 143040 79218
rect 142988 79154 143040 79160
rect 142908 79070 143028 79098
rect 142816 78934 142936 78962
rect 142908 70990 142936 78934
rect 143000 78538 143028 79070
rect 142988 78532 143040 78538
rect 142988 78474 143040 78480
rect 142988 78396 143040 78402
rect 142988 78338 143040 78344
rect 143000 73778 143028 78338
rect 142988 73772 143040 73778
rect 142988 73714 143040 73720
rect 142896 70984 142948 70990
rect 142896 70926 142948 70932
rect 143000 70802 143028 73714
rect 143092 72826 143120 79426
rect 143184 74526 143212 79648
rect 143356 79630 143408 79636
rect 143264 79552 143316 79558
rect 143264 79494 143316 79500
rect 143172 74520 143224 74526
rect 143172 74462 143224 74468
rect 143172 74384 143224 74390
rect 143172 74326 143224 74332
rect 143080 72820 143132 72826
rect 143080 72762 143132 72768
rect 143092 71670 143120 72762
rect 143080 71664 143132 71670
rect 143080 71606 143132 71612
rect 142816 70774 143028 70802
rect 142712 68876 142764 68882
rect 142712 68818 142764 68824
rect 142356 64846 142568 64874
rect 142356 55282 142384 64846
rect 142344 55276 142396 55282
rect 142344 55218 142396 55224
rect 142252 42628 142304 42634
rect 142252 42570 142304 42576
rect 142066 36000 142122 36009
rect 142066 35935 142122 35944
rect 142066 35864 142122 35873
rect 142066 35799 142122 35808
rect 142080 26353 142108 35799
rect 142066 26344 142122 26353
rect 142066 26279 142122 26288
rect 142066 26208 142122 26217
rect 142066 26143 142122 26152
rect 142080 16697 142108 26143
rect 142066 16688 142122 16697
rect 142066 16623 142122 16632
rect 142066 16552 142122 16561
rect 142066 16487 142122 16496
rect 142080 7041 142108 16487
rect 142066 7032 142122 7041
rect 142066 6967 142122 6976
rect 142066 6896 142122 6905
rect 142066 6831 142122 6840
rect 142080 3369 142108 6831
rect 142816 4214 142844 70774
rect 142988 70712 143040 70718
rect 142988 70654 143040 70660
rect 143000 61946 143028 70654
rect 142988 61940 143040 61946
rect 142988 61882 143040 61888
rect 143184 6914 143212 74326
rect 143276 69970 143304 79494
rect 143368 78606 143396 79630
rect 143356 78600 143408 78606
rect 143356 78542 143408 78548
rect 143460 78130 143488 79698
rect 143690 79676 143718 79902
rect 143768 79863 143824 79872
rect 143874 79830 143902 80036
rect 143966 79898 143994 80036
rect 143954 79892 144006 79898
rect 143954 79834 144006 79840
rect 143862 79824 143914 79830
rect 143862 79766 143914 79772
rect 144058 79744 144086 80036
rect 144150 79966 144178 80036
rect 144242 79966 144270 80036
rect 144138 79960 144190 79966
rect 144138 79902 144190 79908
rect 144230 79960 144282 79966
rect 144230 79902 144282 79908
rect 144334 79830 144362 80036
rect 144426 79830 144454 80036
rect 144518 79830 144546 80036
rect 144610 79898 144638 80036
rect 144598 79892 144650 79898
rect 144598 79834 144650 79840
rect 144184 79824 144236 79830
rect 144184 79766 144236 79772
rect 144322 79824 144374 79830
rect 144322 79766 144374 79772
rect 144414 79824 144466 79830
rect 144414 79766 144466 79772
rect 144506 79824 144558 79830
rect 144702 79801 144730 80036
rect 144794 79971 144822 80036
rect 144780 79962 144836 79971
rect 144780 79897 144836 79906
rect 144886 79898 144914 80036
rect 144978 79966 145006 80036
rect 144966 79960 145018 79966
rect 144966 79902 145018 79908
rect 144874 79892 144926 79898
rect 144874 79834 144926 79840
rect 144506 79766 144558 79772
rect 144688 79792 144744 79801
rect 144012 79716 144086 79744
rect 143538 79656 143594 79665
rect 143538 79591 143594 79600
rect 143644 79648 143718 79676
rect 143908 79688 143960 79694
rect 143552 78402 143580 79591
rect 143540 78396 143592 78402
rect 143540 78338 143592 78344
rect 143448 78124 143500 78130
rect 143448 78066 143500 78072
rect 143460 74390 143488 78066
rect 143540 76696 143592 76702
rect 143540 76638 143592 76644
rect 143448 74384 143500 74390
rect 143448 74326 143500 74332
rect 143264 69964 143316 69970
rect 143264 69906 143316 69912
rect 143552 8974 143580 76638
rect 143644 28966 143672 79648
rect 143908 79630 143960 79636
rect 143816 79552 143868 79558
rect 143816 79494 143868 79500
rect 143724 79484 143776 79490
rect 143724 79426 143776 79432
rect 143736 78713 143764 79426
rect 143828 78985 143856 79494
rect 143814 78976 143870 78985
rect 143814 78911 143870 78920
rect 143722 78704 143778 78713
rect 143722 78639 143778 78648
rect 143736 37942 143764 78639
rect 143828 46918 143856 78911
rect 143920 74254 143948 79630
rect 144012 74594 144040 79716
rect 144092 79620 144144 79626
rect 144092 79562 144144 79568
rect 144104 78266 144132 79562
rect 144092 78260 144144 78266
rect 144092 78202 144144 78208
rect 144104 76702 144132 78202
rect 144196 76974 144224 79766
rect 145070 79744 145098 80036
rect 145162 79778 145190 80036
rect 145254 79971 145282 80036
rect 145240 79962 145296 79971
rect 145346 79966 145374 80036
rect 145240 79897 145296 79906
rect 145334 79960 145386 79966
rect 145334 79902 145386 79908
rect 145438 79898 145466 80036
rect 145426 79892 145478 79898
rect 145426 79834 145478 79840
rect 145530 79778 145558 80036
rect 145622 79937 145650 80036
rect 145608 79928 145664 79937
rect 145714 79898 145742 80036
rect 145806 79966 145834 80036
rect 145898 79966 145926 80036
rect 145794 79960 145846 79966
rect 145794 79902 145846 79908
rect 145886 79960 145938 79966
rect 145990 79937 146018 80036
rect 146082 79966 146110 80036
rect 146070 79960 146122 79966
rect 145886 79902 145938 79908
rect 145976 79928 146032 79937
rect 145608 79863 145664 79872
rect 145702 79892 145754 79898
rect 146174 79937 146202 80036
rect 146266 79966 146294 80036
rect 146254 79960 146306 79966
rect 146070 79902 146122 79908
rect 146160 79928 146216 79937
rect 145976 79863 146032 79872
rect 146254 79902 146306 79908
rect 146358 79898 146386 80036
rect 146450 79898 146478 80036
rect 146542 79966 146570 80036
rect 146530 79960 146582 79966
rect 146634 79937 146662 80036
rect 146530 79902 146582 79908
rect 146620 79928 146676 79937
rect 146160 79863 146216 79872
rect 146346 79892 146398 79898
rect 145702 79834 145754 79840
rect 146346 79834 146398 79840
rect 146438 79892 146490 79898
rect 146620 79863 146676 79872
rect 146438 79834 146490 79840
rect 145162 79750 145236 79778
rect 144688 79727 144744 79736
rect 145024 79716 145098 79744
rect 144736 79688 144788 79694
rect 144366 79656 144422 79665
rect 144276 79620 144328 79626
rect 145024 79642 145052 79716
rect 144736 79630 144788 79636
rect 144366 79591 144422 79600
rect 144276 79562 144328 79568
rect 144184 76968 144236 76974
rect 144184 76910 144236 76916
rect 144092 76696 144144 76702
rect 144092 76638 144144 76644
rect 144000 74588 144052 74594
rect 144000 74530 144052 74536
rect 143908 74248 143960 74254
rect 143908 74190 143960 74196
rect 144012 72962 144040 74530
rect 144288 74474 144316 79562
rect 144380 74534 144408 79591
rect 144644 79552 144696 79558
rect 144644 79494 144696 79500
rect 144552 79484 144604 79490
rect 144552 79426 144604 79432
rect 144460 77172 144512 77178
rect 144460 77114 144512 77120
rect 144472 75886 144500 77114
rect 144460 75880 144512 75886
rect 144460 75822 144512 75828
rect 144564 74769 144592 79426
rect 144550 74760 144606 74769
rect 144550 74695 144606 74704
rect 144380 74506 144592 74534
rect 144104 74446 144316 74474
rect 144104 73166 144132 74446
rect 144564 74186 144592 74506
rect 144656 74458 144684 79494
rect 144748 75177 144776 79630
rect 144828 79620 144880 79626
rect 144828 79562 144880 79568
rect 144932 79614 145052 79642
rect 144840 79257 144868 79562
rect 144826 79248 144882 79257
rect 144826 79183 144882 79192
rect 144734 75168 144790 75177
rect 144734 75103 144790 75112
rect 144644 74452 144696 74458
rect 144644 74394 144696 74400
rect 144552 74180 144604 74186
rect 144552 74122 144604 74128
rect 144092 73160 144144 73166
rect 144092 73102 144144 73108
rect 144000 72956 144052 72962
rect 144000 72898 144052 72904
rect 144104 71774 144132 73102
rect 144276 72956 144328 72962
rect 144276 72898 144328 72904
rect 144012 71746 144132 71774
rect 144012 66230 144040 71746
rect 144288 70854 144316 72898
rect 144276 70848 144328 70854
rect 144276 70790 144328 70796
rect 144564 70106 144592 74122
rect 144552 70100 144604 70106
rect 144552 70042 144604 70048
rect 144000 66224 144052 66230
rect 144000 66166 144052 66172
rect 144656 61538 144684 74394
rect 144748 71097 144776 75103
rect 144734 71088 144790 71097
rect 144734 71023 144790 71032
rect 144644 61532 144696 61538
rect 144644 61474 144696 61480
rect 144840 57974 144868 79183
rect 144932 74322 144960 79614
rect 145208 75478 145236 79750
rect 145392 79750 145558 79778
rect 145746 79792 145802 79801
rect 145930 79792 145986 79801
rect 145392 78946 145420 79750
rect 145746 79727 145748 79736
rect 145800 79727 145802 79736
rect 145840 79756 145892 79762
rect 145748 79698 145800 79704
rect 145930 79727 145986 79736
rect 146114 79792 146170 79801
rect 146726 79778 146754 80036
rect 146818 79966 146846 80036
rect 146910 79971 146938 80172
rect 177764 80096 177816 80102
rect 177764 80038 177816 80044
rect 146806 79960 146858 79966
rect 146806 79902 146858 79908
rect 146896 79962 146952 79971
rect 147002 79966 147030 80036
rect 147094 79966 147122 80036
rect 147186 79966 147214 80036
rect 146896 79897 146952 79906
rect 146990 79960 147042 79966
rect 146990 79902 147042 79908
rect 147082 79960 147134 79966
rect 147082 79902 147134 79908
rect 147174 79960 147226 79966
rect 147278 79937 147306 80036
rect 147370 79966 147398 80036
rect 147358 79960 147410 79966
rect 147174 79902 147226 79908
rect 147264 79928 147320 79937
rect 147358 79902 147410 79908
rect 147462 79898 147490 80036
rect 147264 79863 147320 79872
rect 147450 79892 147502 79898
rect 147450 79834 147502 79840
rect 147036 79824 147088 79830
rect 146942 79792 146998 79801
rect 146170 79750 146248 79778
rect 146114 79727 146170 79736
rect 145840 79698 145892 79704
rect 145472 79688 145524 79694
rect 145656 79688 145708 79694
rect 145524 79648 145604 79676
rect 145472 79630 145524 79636
rect 145380 78940 145432 78946
rect 145380 78882 145432 78888
rect 145196 75472 145248 75478
rect 145196 75414 145248 75420
rect 145104 75336 145156 75342
rect 145104 75278 145156 75284
rect 144920 74316 144972 74322
rect 144920 74258 144972 74264
rect 144932 67590 144960 74258
rect 145012 72412 145064 72418
rect 145012 72354 145064 72360
rect 144920 67584 144972 67590
rect 144920 67526 144972 67532
rect 144840 57946 144960 57974
rect 143816 46912 143868 46918
rect 143816 46854 143868 46860
rect 143724 37936 143776 37942
rect 143724 37878 143776 37884
rect 144932 35222 144960 57946
rect 145024 47598 145052 72354
rect 145116 51882 145144 75278
rect 145208 60178 145236 75414
rect 145392 72418 145420 78882
rect 145576 75206 145604 79648
rect 145656 79630 145708 79636
rect 145668 77178 145696 79630
rect 145656 77172 145708 77178
rect 145656 77114 145708 77120
rect 145760 75342 145788 79698
rect 145748 75336 145800 75342
rect 145748 75278 145800 75284
rect 145564 75200 145616 75206
rect 145564 75142 145616 75148
rect 145380 72412 145432 72418
rect 145380 72354 145432 72360
rect 145196 60172 145248 60178
rect 145196 60114 145248 60120
rect 145104 51876 145156 51882
rect 145104 51818 145156 51824
rect 145012 47592 145064 47598
rect 145012 47534 145064 47540
rect 144920 35216 144972 35222
rect 144920 35158 144972 35164
rect 143632 28960 143684 28966
rect 143632 28902 143684 28908
rect 144920 28960 144972 28966
rect 144920 28902 144972 28908
rect 144932 16574 144960 28902
rect 145576 17270 145604 75142
rect 145852 73953 145880 79698
rect 145944 75449 145972 79727
rect 146024 79688 146076 79694
rect 146024 79630 146076 79636
rect 146116 79688 146168 79694
rect 146116 79630 146168 79636
rect 146036 77450 146064 79630
rect 146024 77444 146076 77450
rect 146024 77386 146076 77392
rect 146036 75954 146064 77386
rect 146024 75948 146076 75954
rect 146024 75890 146076 75896
rect 145930 75440 145986 75449
rect 145930 75375 145986 75384
rect 146128 75313 146156 79630
rect 146114 75304 146170 75313
rect 146114 75239 146170 75248
rect 145838 73944 145894 73953
rect 145838 73879 145894 73888
rect 146220 24138 146248 79750
rect 146300 79756 146352 79762
rect 146300 79698 146352 79704
rect 146392 79756 146444 79762
rect 146392 79698 146444 79704
rect 146576 79756 146628 79762
rect 146726 79750 146800 79778
rect 146576 79698 146628 79704
rect 146312 78674 146340 79698
rect 146300 78668 146352 78674
rect 146300 78610 146352 78616
rect 146404 75750 146432 79698
rect 146482 79656 146538 79665
rect 146482 79591 146538 79600
rect 146392 75744 146444 75750
rect 146392 75686 146444 75692
rect 146300 70100 146352 70106
rect 146300 70042 146352 70048
rect 146208 24132 146260 24138
rect 146208 24074 146260 24080
rect 145564 17264 145616 17270
rect 145564 17206 145616 17212
rect 146312 16574 146340 70042
rect 146496 65550 146524 79591
rect 146588 75546 146616 79698
rect 146668 79688 146720 79694
rect 146668 79630 146720 79636
rect 146680 76430 146708 79630
rect 146772 78577 146800 79750
rect 147036 79766 147088 79772
rect 147220 79824 147272 79830
rect 147220 79766 147272 79772
rect 147312 79824 147364 79830
rect 147312 79766 147364 79772
rect 146942 79727 146998 79736
rect 146852 79688 146904 79694
rect 146852 79630 146904 79636
rect 146864 78742 146892 79630
rect 146852 78736 146904 78742
rect 146852 78678 146904 78684
rect 146758 78568 146814 78577
rect 146758 78503 146814 78512
rect 146668 76424 146720 76430
rect 146668 76366 146720 76372
rect 146772 75682 146800 78503
rect 146956 77625 146984 79727
rect 146942 77616 146998 77625
rect 146942 77551 146998 77560
rect 146944 75948 146996 75954
rect 146944 75890 146996 75896
rect 146760 75676 146812 75682
rect 146760 75618 146812 75624
rect 146576 75540 146628 75546
rect 146576 75482 146628 75488
rect 146484 65544 146536 65550
rect 146484 65486 146536 65492
rect 144932 16546 145512 16574
rect 146312 16546 146892 16574
rect 143540 8968 143592 8974
rect 143540 8910 143592 8916
rect 142908 6886 143212 6914
rect 142804 4208 142856 4214
rect 142804 4150 142856 4156
rect 142908 3482 142936 6886
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 142448 3454 142936 3482
rect 142066 3360 142122 3369
rect 142066 3295 142122 3304
rect 141424 3052 141476 3058
rect 141424 2994 141476 3000
rect 140792 1278 141280 1306
rect 141252 480 141280 1278
rect 142448 480 142476 3454
rect 143552 480 143580 4150
rect 144736 4004 144788 4010
rect 144736 3946 144788 3952
rect 144748 480 144776 3946
rect 140014 354 140126 480
rect 139412 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 146864 3482 146892 16546
rect 146956 4146 146984 75890
rect 147048 74338 147076 79766
rect 147128 79484 147180 79490
rect 147128 79426 147180 79432
rect 147140 79257 147168 79426
rect 147126 79248 147182 79257
rect 147126 79183 147182 79192
rect 147232 79082 147260 79766
rect 147220 79076 147272 79082
rect 147220 79018 147272 79024
rect 147232 78606 147260 79018
rect 147220 78600 147272 78606
rect 147220 78542 147272 78548
rect 147324 76945 147352 79766
rect 147404 79756 147456 79762
rect 147554 79744 147582 80036
rect 147404 79698 147456 79704
rect 147508 79716 147582 79744
rect 147646 79744 147674 80036
rect 147738 79812 147766 80036
rect 147830 79966 147858 80036
rect 147818 79960 147870 79966
rect 147818 79902 147870 79908
rect 147738 79784 147812 79812
rect 147646 79716 147720 79744
rect 147416 79150 147444 79698
rect 147404 79144 147456 79150
rect 147508 79121 147536 79716
rect 147586 79656 147642 79665
rect 147586 79591 147642 79600
rect 147404 79086 147456 79092
rect 147494 79112 147550 79121
rect 147310 76936 147366 76945
rect 147310 76871 147366 76880
rect 147048 74310 147260 74338
rect 147128 74248 147180 74254
rect 147128 74190 147180 74196
rect 147140 70938 147168 74190
rect 147048 70910 147168 70938
rect 146944 4140 146996 4146
rect 146944 4082 146996 4088
rect 147048 3670 147076 70910
rect 147128 70848 147180 70854
rect 147128 70790 147180 70796
rect 147140 3738 147168 70790
rect 147232 70009 147260 74310
rect 147218 70000 147274 70009
rect 147218 69935 147274 69944
rect 147220 67584 147272 67590
rect 147220 67526 147272 67532
rect 147232 3806 147260 67526
rect 147312 60172 147364 60178
rect 147312 60114 147364 60120
rect 147324 4078 147352 60114
rect 147416 58750 147444 79086
rect 147494 79047 147550 79056
rect 147404 58744 147456 58750
rect 147404 58686 147456 58692
rect 147600 51746 147628 79591
rect 147692 77081 147720 79716
rect 147784 79506 147812 79784
rect 147922 79778 147950 80036
rect 148014 79966 148042 80036
rect 148106 79966 148134 80036
rect 148198 79966 148226 80036
rect 148002 79960 148054 79966
rect 148002 79902 148054 79908
rect 148094 79960 148146 79966
rect 148094 79902 148146 79908
rect 148186 79960 148238 79966
rect 148186 79902 148238 79908
rect 148290 79898 148318 80036
rect 148382 79898 148410 80036
rect 148474 79971 148502 80036
rect 148460 79962 148516 79971
rect 148278 79892 148330 79898
rect 148278 79834 148330 79840
rect 148370 79892 148422 79898
rect 148460 79897 148516 79906
rect 148566 79898 148594 80036
rect 148658 79971 148686 80036
rect 148644 79962 148700 79971
rect 148750 79966 148778 80036
rect 148370 79834 148422 79840
rect 148554 79892 148606 79898
rect 148644 79897 148700 79906
rect 148738 79960 148790 79966
rect 148738 79902 148790 79908
rect 148842 79898 148870 80036
rect 148934 79937 148962 80036
rect 148920 79928 148976 79937
rect 148554 79834 148606 79840
rect 148830 79892 148882 79898
rect 148920 79863 148976 79872
rect 148830 79834 148882 79840
rect 148692 79824 148744 79830
rect 147876 79750 147950 79778
rect 148046 79792 148102 79801
rect 147876 79626 147904 79750
rect 148046 79727 148048 79736
rect 148100 79727 148102 79736
rect 148230 79792 148286 79801
rect 148286 79750 148456 79778
rect 148744 79772 148824 79778
rect 148692 79766 148824 79772
rect 148230 79727 148286 79736
rect 148048 79698 148100 79704
rect 147956 79688 148008 79694
rect 147956 79630 148008 79636
rect 147864 79620 147916 79626
rect 147864 79562 147916 79568
rect 147784 79478 147904 79506
rect 147876 79014 147904 79478
rect 147968 79286 147996 79630
rect 147956 79280 148008 79286
rect 147956 79222 148008 79228
rect 147864 79008 147916 79014
rect 147864 78950 147916 78956
rect 147772 77104 147824 77110
rect 147678 77072 147734 77081
rect 147772 77046 147824 77052
rect 147678 77007 147734 77016
rect 147588 51740 147640 51746
rect 147588 51682 147640 51688
rect 147784 47802 147812 77046
rect 147876 55962 147904 78950
rect 147968 77110 147996 79222
rect 147956 77104 148008 77110
rect 147956 77046 148008 77052
rect 148060 75546 148088 79698
rect 148140 79688 148192 79694
rect 148140 79630 148192 79636
rect 148324 79688 148376 79694
rect 148324 79630 148376 79636
rect 148152 75993 148180 79630
rect 148336 78198 148364 79630
rect 148324 78192 148376 78198
rect 148324 78134 148376 78140
rect 148336 76702 148364 78134
rect 148428 77926 148456 79750
rect 148600 79756 148652 79762
rect 148704 79750 148824 79766
rect 148600 79698 148652 79704
rect 148508 79552 148560 79558
rect 148508 79494 148560 79500
rect 148520 78334 148548 79494
rect 148508 78328 148560 78334
rect 148508 78270 148560 78276
rect 148416 77920 148468 77926
rect 148416 77862 148468 77868
rect 148414 77752 148470 77761
rect 148414 77687 148470 77696
rect 148324 76696 148376 76702
rect 148324 76638 148376 76644
rect 148138 75984 148194 75993
rect 148138 75919 148194 75928
rect 147956 75540 148008 75546
rect 147956 75482 148008 75488
rect 148048 75540 148100 75546
rect 148048 75482 148100 75488
rect 147968 69698 147996 75482
rect 148428 70394 148456 77687
rect 148152 70366 148456 70394
rect 147956 69692 148008 69698
rect 147956 69634 148008 69640
rect 147864 55956 147916 55962
rect 147864 55898 147916 55904
rect 148152 54602 148180 70366
rect 148322 68912 148378 68921
rect 148322 68847 148378 68856
rect 148140 54596 148192 54602
rect 148140 54538 148192 54544
rect 147772 47796 147824 47802
rect 147772 47738 147824 47744
rect 147772 46912 147824 46918
rect 147772 46854 147824 46860
rect 147784 16574 147812 46854
rect 147784 16546 147904 16574
rect 147404 4140 147456 4146
rect 147404 4082 147456 4088
rect 147312 4072 147364 4078
rect 147312 4014 147364 4020
rect 147220 3800 147272 3806
rect 147220 3742 147272 3748
rect 147128 3732 147180 3738
rect 147128 3674 147180 3680
rect 147036 3664 147088 3670
rect 147036 3606 147088 3612
rect 146864 3454 147168 3482
rect 147140 480 147168 3454
rect 147416 3398 147444 4082
rect 147404 3392 147456 3398
rect 147404 3334 147456 3340
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 148336 3466 148364 68847
rect 148416 66224 148468 66230
rect 148416 66166 148468 66172
rect 148324 3460 148376 3466
rect 148324 3402 148376 3408
rect 148428 3194 148456 66166
rect 148520 41002 148548 78270
rect 148612 76770 148640 79698
rect 148692 79620 148744 79626
rect 148692 79562 148744 79568
rect 148704 78946 148732 79562
rect 148692 78940 148744 78946
rect 148692 78882 148744 78888
rect 148796 78305 148824 79750
rect 149026 79744 149054 80036
rect 149118 79937 149146 80036
rect 149210 79966 149238 80036
rect 149198 79960 149250 79966
rect 149104 79928 149160 79937
rect 149198 79902 149250 79908
rect 149302 79898 149330 80036
rect 149394 79898 149422 80036
rect 149104 79863 149160 79872
rect 149290 79892 149342 79898
rect 149290 79834 149342 79840
rect 149382 79892 149434 79898
rect 149382 79834 149434 79840
rect 148980 79716 149054 79744
rect 149244 79756 149296 79762
rect 148876 79484 148928 79490
rect 148876 79426 148928 79432
rect 148782 78296 148838 78305
rect 148782 78231 148838 78240
rect 148784 77920 148836 77926
rect 148784 77862 148836 77868
rect 148796 76838 148824 77862
rect 148784 76832 148836 76838
rect 148784 76774 148836 76780
rect 148600 76764 148652 76770
rect 148600 76706 148652 76712
rect 148612 47734 148640 76706
rect 148692 76696 148744 76702
rect 148692 76638 148744 76644
rect 148704 55894 148732 76638
rect 148796 65618 148824 76774
rect 148784 65612 148836 65618
rect 148784 65554 148836 65560
rect 148692 55888 148744 55894
rect 148692 55830 148744 55836
rect 148600 47728 148652 47734
rect 148600 47670 148652 47676
rect 148508 40996 148560 41002
rect 148508 40938 148560 40944
rect 148888 31414 148916 79426
rect 148980 79121 149008 79716
rect 149486 79744 149514 80036
rect 149296 79716 149376 79744
rect 149244 79698 149296 79704
rect 149242 79656 149298 79665
rect 149242 79591 149298 79600
rect 149256 79354 149284 79591
rect 149244 79348 149296 79354
rect 149244 79290 149296 79296
rect 148966 79112 149022 79121
rect 148966 79047 149022 79056
rect 149150 79112 149206 79121
rect 149150 79047 149206 79056
rect 149060 78804 149112 78810
rect 149060 78746 149112 78752
rect 148968 78668 149020 78674
rect 148968 78610 149020 78616
rect 148980 71126 149008 78610
rect 148968 71120 149020 71126
rect 148968 71062 149020 71068
rect 149072 36786 149100 78746
rect 149060 36780 149112 36786
rect 149060 36722 149112 36728
rect 148876 31408 148928 31414
rect 148876 31350 148928 31356
rect 149164 7818 149192 79047
rect 149256 53242 149284 79290
rect 149348 76702 149376 79716
rect 149440 79716 149514 79744
rect 149440 77897 149468 79716
rect 149578 79676 149606 80036
rect 149670 79744 149698 80036
rect 149762 79812 149790 80036
rect 149854 79966 149882 80036
rect 149842 79960 149894 79966
rect 149842 79902 149894 79908
rect 149946 79812 149974 80036
rect 150038 79898 150066 80036
rect 150130 79966 150158 80036
rect 150118 79960 150170 79966
rect 150222 79937 150250 80036
rect 150314 79966 150342 80036
rect 150302 79960 150354 79966
rect 150118 79902 150170 79908
rect 150208 79928 150264 79937
rect 150026 79892 150078 79898
rect 150406 79937 150434 80036
rect 150302 79902 150354 79908
rect 150392 79928 150448 79937
rect 150208 79863 150264 79872
rect 150392 79863 150448 79872
rect 150026 79834 150078 79840
rect 149762 79784 149836 79812
rect 149670 79716 149744 79744
rect 149532 79648 149606 79676
rect 149716 79665 149744 79716
rect 149702 79656 149758 79665
rect 149426 77888 149482 77897
rect 149426 77823 149482 77832
rect 149440 76906 149468 77823
rect 149428 76900 149480 76906
rect 149428 76842 149480 76848
rect 149336 76696 149388 76702
rect 149336 76638 149388 76644
rect 149336 73092 149388 73098
rect 149336 73034 149388 73040
rect 149348 64874 149376 73034
rect 149532 72554 149560 79648
rect 149702 79591 149758 79600
rect 149716 79506 149744 79591
rect 149624 79478 149744 79506
rect 149624 76634 149652 79478
rect 149704 79416 149756 79422
rect 149704 79358 149756 79364
rect 149716 78130 149744 79358
rect 149704 78124 149756 78130
rect 149704 78066 149756 78072
rect 149612 76628 149664 76634
rect 149612 76570 149664 76576
rect 149520 72548 149572 72554
rect 149520 72490 149572 72496
rect 149808 71534 149836 79784
rect 149900 79784 149974 79812
rect 150256 79824 150308 79830
rect 150254 79792 150256 79801
rect 150308 79792 150310 79801
rect 149900 79608 149928 79784
rect 150254 79727 150310 79736
rect 150348 79756 150400 79762
rect 150498 79744 150526 80036
rect 150348 79698 150400 79704
rect 150452 79716 150526 79744
rect 150590 79744 150618 80036
rect 150682 79966 150710 80036
rect 150670 79960 150722 79966
rect 150670 79902 150722 79908
rect 150774 79744 150802 80036
rect 150866 79971 150894 80036
rect 150852 79962 150908 79971
rect 150958 79966 150986 80036
rect 150852 79897 150908 79906
rect 150946 79960 150998 79966
rect 150946 79902 150998 79908
rect 151050 79801 151078 80036
rect 151142 79937 151170 80036
rect 151128 79928 151184 79937
rect 151128 79863 151130 79872
rect 151182 79863 151184 79872
rect 151130 79834 151182 79840
rect 151142 79803 151170 79834
rect 150898 79792 150954 79801
rect 150590 79716 150664 79744
rect 150774 79716 150848 79744
rect 150898 79727 150954 79736
rect 151036 79792 151092 79801
rect 151234 79744 151262 80036
rect 151326 79830 151354 80036
rect 151418 79966 151446 80036
rect 151406 79960 151458 79966
rect 151406 79902 151458 79908
rect 151510 79898 151538 80036
rect 151498 79892 151550 79898
rect 151498 79834 151550 79840
rect 151314 79824 151366 79830
rect 151314 79766 151366 79772
rect 151036 79727 151092 79736
rect 150164 79688 150216 79694
rect 150164 79630 150216 79636
rect 149900 79580 150112 79608
rect 149980 79484 150032 79490
rect 149980 79426 150032 79432
rect 149888 79416 149940 79422
rect 149888 79358 149940 79364
rect 149900 73098 149928 79358
rect 149992 78690 150020 79426
rect 150084 78810 150112 79580
rect 150072 78804 150124 78810
rect 150072 78746 150124 78752
rect 149992 78662 150112 78690
rect 150084 78169 150112 78662
rect 150176 78305 150204 79630
rect 150162 78296 150218 78305
rect 150162 78231 150218 78240
rect 150070 78160 150126 78169
rect 150070 78095 150126 78104
rect 149980 76900 150032 76906
rect 149980 76842 150032 76848
rect 149888 73092 149940 73098
rect 149888 73034 149940 73040
rect 149888 72548 149940 72554
rect 149888 72490 149940 72496
rect 149796 71528 149848 71534
rect 149796 71470 149848 71476
rect 149348 64846 149744 64874
rect 149716 64326 149744 64846
rect 149704 64320 149756 64326
rect 149704 64262 149756 64268
rect 149704 61532 149756 61538
rect 149704 61474 149756 61480
rect 149244 53236 149296 53242
rect 149244 53178 149296 53184
rect 149152 7812 149204 7818
rect 149152 7754 149204 7760
rect 149716 4010 149744 61474
rect 149808 60246 149836 71470
rect 149900 68474 149928 72490
rect 149888 68468 149940 68474
rect 149888 68410 149940 68416
rect 149796 60240 149848 60246
rect 149796 60182 149848 60188
rect 149794 50688 149850 50697
rect 149794 50623 149850 50632
rect 149704 4004 149756 4010
rect 149704 3946 149756 3952
rect 149808 3942 149836 50623
rect 149992 23050 150020 76842
rect 150084 70394 150112 78095
rect 150256 76628 150308 76634
rect 150256 76570 150308 76576
rect 150084 70366 150204 70394
rect 150176 50522 150204 70366
rect 150164 50516 150216 50522
rect 150164 50458 150216 50464
rect 150268 49162 150296 76570
rect 150360 75478 150388 79698
rect 150452 77858 150480 79716
rect 150530 79656 150586 79665
rect 150530 79591 150532 79600
rect 150584 79591 150586 79600
rect 150532 79562 150584 79568
rect 150532 78600 150584 78606
rect 150532 78542 150584 78548
rect 150440 77852 150492 77858
rect 150440 77794 150492 77800
rect 150348 75472 150400 75478
rect 150348 75414 150400 75420
rect 150544 64190 150572 78542
rect 150636 78266 150664 79716
rect 150716 79620 150768 79626
rect 150716 79562 150768 79568
rect 150624 78260 150676 78266
rect 150624 78202 150676 78208
rect 150728 70394 150756 79562
rect 150820 79490 150848 79716
rect 150912 79676 150940 79727
rect 151188 79716 151262 79744
rect 151452 79756 151504 79762
rect 150912 79648 151032 79676
rect 150900 79552 150952 79558
rect 150900 79494 150952 79500
rect 150808 79484 150860 79490
rect 150808 79426 150860 79432
rect 150806 79384 150862 79393
rect 150806 79319 150862 79328
rect 150636 70366 150756 70394
rect 150532 64184 150584 64190
rect 150532 64126 150584 64132
rect 150256 49156 150308 49162
rect 150256 49098 150308 49104
rect 149980 23044 150032 23050
rect 149980 22986 150032 22992
rect 150636 17542 150664 70366
rect 150820 60178 150848 79319
rect 150808 60172 150860 60178
rect 150808 60114 150860 60120
rect 150624 17536 150676 17542
rect 150624 17478 150676 17484
rect 150912 11966 150940 79494
rect 151004 74254 151032 79648
rect 151082 79656 151138 79665
rect 151082 79591 151138 79600
rect 151096 78418 151124 79591
rect 151188 78713 151216 79716
rect 151602 79744 151630 80036
rect 151694 79971 151722 80036
rect 151680 79962 151736 79971
rect 151680 79897 151736 79906
rect 151786 79778 151814 80036
rect 151878 79971 151906 80036
rect 151864 79962 151920 79971
rect 151864 79897 151920 79906
rect 151740 79750 151814 79778
rect 151602 79716 151676 79744
rect 151452 79698 151504 79704
rect 151360 79688 151412 79694
rect 151266 79656 151322 79665
rect 151360 79630 151412 79636
rect 151266 79591 151268 79600
rect 151320 79591 151322 79600
rect 151268 79562 151320 79568
rect 151174 78704 151230 78713
rect 151174 78639 151230 78648
rect 151096 78390 151308 78418
rect 151176 78260 151228 78266
rect 151176 78202 151228 78208
rect 151084 75880 151136 75886
rect 151084 75822 151136 75828
rect 150992 74248 151044 74254
rect 150992 74190 151044 74196
rect 150900 11960 150952 11966
rect 150900 11902 150952 11908
rect 150716 4072 150768 4078
rect 150716 4014 150768 4020
rect 149796 3936 149848 3942
rect 149796 3878 149848 3884
rect 150728 3738 150756 4014
rect 150624 3732 150676 3738
rect 150624 3674 150676 3680
rect 150716 3732 150768 3738
rect 150716 3674 150768 3680
rect 149520 3664 149572 3670
rect 149520 3606 149572 3612
rect 148416 3188 148468 3194
rect 148416 3130 148468 3136
rect 149532 480 149560 3606
rect 150636 480 150664 3674
rect 151096 3670 151124 75822
rect 151188 68950 151216 78202
rect 151280 76566 151308 78390
rect 151268 76560 151320 76566
rect 151268 76502 151320 76508
rect 151372 73930 151400 79630
rect 151464 79393 151492 79698
rect 151544 79484 151596 79490
rect 151544 79426 151596 79432
rect 151450 79384 151506 79393
rect 151450 79319 151506 79328
rect 151452 79280 151504 79286
rect 151452 79222 151504 79228
rect 151464 78169 151492 79222
rect 151450 78160 151506 78169
rect 151450 78095 151506 78104
rect 151452 77852 151504 77858
rect 151452 77794 151504 77800
rect 151280 73902 151400 73930
rect 151280 71262 151308 73902
rect 151360 71664 151412 71670
rect 151360 71606 151412 71612
rect 151268 71256 151320 71262
rect 151268 71198 151320 71204
rect 151176 68944 151228 68950
rect 151176 68886 151228 68892
rect 151188 9314 151216 68886
rect 151280 28558 151308 71198
rect 151372 71194 151400 71606
rect 151360 71188 151412 71194
rect 151360 71130 151412 71136
rect 151372 46442 151400 71130
rect 151464 57322 151492 77794
rect 151556 71670 151584 79426
rect 151648 76401 151676 79716
rect 151740 79490 151768 79750
rect 151970 79744 151998 80036
rect 152062 79966 152090 80036
rect 152050 79960 152102 79966
rect 152050 79902 152102 79908
rect 152154 79744 152182 80036
rect 152246 79801 152274 80036
rect 151970 79716 152044 79744
rect 151910 79656 151966 79665
rect 151910 79591 151966 79600
rect 151728 79484 151780 79490
rect 151728 79426 151780 79432
rect 151726 78432 151782 78441
rect 151726 78367 151782 78376
rect 151634 76392 151690 76401
rect 151634 76327 151690 76336
rect 151740 73846 151768 78367
rect 151820 76968 151872 76974
rect 151820 76910 151872 76916
rect 151728 73840 151780 73846
rect 151728 73782 151780 73788
rect 151544 71664 151596 71670
rect 151544 71606 151596 71612
rect 151452 57316 151504 57322
rect 151452 57258 151504 57264
rect 151360 46436 151412 46442
rect 151360 46378 151412 46384
rect 151268 28552 151320 28558
rect 151268 28494 151320 28500
rect 151176 9308 151228 9314
rect 151176 9250 151228 9256
rect 151832 4078 151860 76910
rect 151924 71738 151952 79591
rect 152016 78810 152044 79716
rect 152108 79716 152182 79744
rect 152232 79792 152288 79801
rect 152232 79727 152288 79736
rect 152108 79490 152136 79716
rect 152338 79676 152366 80036
rect 152430 79744 152458 80036
rect 152522 79903 152550 80036
rect 152508 79894 152564 79903
rect 152508 79829 152564 79838
rect 152614 79778 152642 80036
rect 152706 79898 152734 80036
rect 152694 79892 152746 79898
rect 152694 79834 152746 79840
rect 152798 79778 152826 80036
rect 152568 79750 152642 79778
rect 152752 79750 152826 79778
rect 152430 79716 152504 79744
rect 152338 79648 152412 79676
rect 152280 79552 152332 79558
rect 152280 79494 152332 79500
rect 152096 79484 152148 79490
rect 152096 79426 152148 79432
rect 152186 79384 152242 79393
rect 152108 79328 152186 79336
rect 152108 79308 152188 79328
rect 152004 78804 152056 78810
rect 152004 78746 152056 78752
rect 152004 78668 152056 78674
rect 152004 78610 152056 78616
rect 152016 73030 152044 78610
rect 152004 73024 152056 73030
rect 152004 72966 152056 72972
rect 152016 72282 152044 72966
rect 152004 72276 152056 72282
rect 152004 72218 152056 72224
rect 151912 71732 151964 71738
rect 151912 71674 151964 71680
rect 151924 71194 151952 71674
rect 151912 71188 151964 71194
rect 151912 71130 151964 71136
rect 151912 8968 151964 8974
rect 151912 8910 151964 8916
rect 151820 4072 151872 4078
rect 151820 4014 151872 4020
rect 151084 3664 151136 3670
rect 151084 3606 151136 3612
rect 151924 3482 151952 8910
rect 152108 5030 152136 79308
rect 152240 79319 152242 79328
rect 152188 79290 152240 79296
rect 152188 78804 152240 78810
rect 152188 78746 152240 78752
rect 152200 70394 152228 78746
rect 152292 74497 152320 79494
rect 152384 78674 152412 79648
rect 152372 78668 152424 78674
rect 152372 78610 152424 78616
rect 152370 78568 152426 78577
rect 152370 78503 152426 78512
rect 152278 74488 152334 74497
rect 152278 74423 152334 74432
rect 152292 73681 152320 74423
rect 152384 74186 152412 78503
rect 152372 74180 152424 74186
rect 152372 74122 152424 74128
rect 152278 73672 152334 73681
rect 152278 73607 152334 73616
rect 152476 71398 152504 79716
rect 152568 79626 152596 79750
rect 152646 79656 152702 79665
rect 152556 79620 152608 79626
rect 152646 79591 152702 79600
rect 152556 79562 152608 79568
rect 152660 79506 152688 79591
rect 152752 79529 152780 79750
rect 152890 79608 152918 80036
rect 152982 79676 153010 80036
rect 153074 79966 153102 80036
rect 153166 79966 153194 80036
rect 153258 79966 153286 80036
rect 153062 79960 153114 79966
rect 153062 79902 153114 79908
rect 153154 79960 153206 79966
rect 153154 79902 153206 79908
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 153108 79824 153160 79830
rect 153108 79766 153160 79772
rect 152982 79648 153056 79676
rect 152890 79580 152964 79608
rect 152568 79478 152688 79506
rect 152738 79520 152794 79529
rect 152568 78198 152596 79478
rect 152738 79455 152794 79464
rect 152832 79484 152884 79490
rect 152648 79416 152700 79422
rect 152648 79358 152700 79364
rect 152556 78192 152608 78198
rect 152556 78134 152608 78140
rect 152660 77042 152688 79358
rect 152648 77036 152700 77042
rect 152648 76978 152700 76984
rect 152752 73914 152780 79455
rect 152832 79426 152884 79432
rect 152844 76265 152872 79426
rect 152936 77897 152964 79580
rect 153028 78305 153056 79648
rect 153014 78296 153070 78305
rect 153014 78231 153070 78240
rect 153016 78192 153068 78198
rect 153120 78169 153148 79766
rect 153200 79756 153252 79762
rect 153350 79744 153378 80036
rect 153442 79966 153470 80036
rect 153430 79960 153482 79966
rect 153430 79902 153482 79908
rect 153534 79778 153562 80036
rect 153488 79750 153562 79778
rect 153350 79716 153424 79744
rect 153200 79698 153252 79704
rect 153016 78134 153068 78140
rect 153106 78160 153162 78169
rect 152922 77888 152978 77897
rect 152922 77823 152978 77832
rect 152830 76256 152886 76265
rect 152830 76191 152886 76200
rect 152740 73908 152792 73914
rect 152740 73850 152792 73856
rect 152738 73672 152794 73681
rect 152738 73607 152794 73616
rect 152464 71392 152516 71398
rect 152464 71334 152516 71340
rect 152200 70366 152320 70394
rect 152292 69018 152320 70366
rect 152280 69012 152332 69018
rect 152280 68954 152332 68960
rect 152476 10606 152504 71334
rect 152648 71188 152700 71194
rect 152648 71130 152700 71136
rect 152556 69012 152608 69018
rect 152556 68954 152608 68960
rect 152568 34066 152596 68954
rect 152660 39642 152688 71130
rect 152752 50454 152780 73607
rect 152832 72276 152884 72282
rect 152832 72218 152884 72224
rect 152844 64258 152872 72218
rect 152832 64252 152884 64258
rect 152832 64194 152884 64200
rect 152740 50448 152792 50454
rect 152740 50390 152792 50396
rect 152648 39636 152700 39642
rect 152648 39578 152700 39584
rect 152556 34060 152608 34066
rect 152556 34002 152608 34008
rect 153028 16182 153056 78134
rect 153106 78095 153162 78104
rect 153212 77994 153240 79698
rect 153292 78668 153344 78674
rect 153292 78610 153344 78616
rect 153200 77988 153252 77994
rect 153200 77930 153252 77936
rect 153106 77616 153162 77625
rect 153106 77551 153162 77560
rect 153120 60042 153148 77551
rect 153200 75268 153252 75274
rect 153200 75210 153252 75216
rect 153212 70378 153240 75210
rect 153304 74526 153332 78610
rect 153292 74520 153344 74526
rect 153292 74462 153344 74468
rect 153304 74050 153332 74462
rect 153396 74458 153424 79716
rect 153488 79608 153516 79750
rect 153626 79744 153654 80036
rect 153718 79898 153746 80036
rect 153706 79892 153758 79898
rect 153706 79834 153758 79840
rect 153810 79812 153838 80036
rect 153902 79937 153930 80036
rect 153888 79928 153944 79937
rect 153888 79863 153944 79872
rect 153810 79784 153884 79812
rect 153626 79716 153792 79744
rect 153764 79665 153792 79716
rect 153750 79656 153806 79665
rect 153488 79580 153608 79608
rect 153750 79591 153806 79600
rect 153474 79520 153530 79529
rect 153474 79455 153530 79464
rect 153384 74452 153436 74458
rect 153384 74394 153436 74400
rect 153488 74118 153516 79455
rect 153476 74112 153528 74118
rect 153476 74054 153528 74060
rect 153292 74044 153344 74050
rect 153292 73986 153344 73992
rect 153200 70372 153252 70378
rect 153200 70314 153252 70320
rect 153580 70038 153608 79580
rect 153764 78470 153792 79591
rect 153752 78464 153804 78470
rect 153752 78406 153804 78412
rect 153660 77988 153712 77994
rect 153660 77930 153712 77936
rect 153672 70242 153700 77930
rect 153856 75274 153884 79784
rect 153994 79778 154022 80036
rect 154086 79898 154114 80036
rect 154178 79898 154206 80036
rect 154074 79892 154126 79898
rect 154074 79834 154126 79840
rect 154166 79892 154218 79898
rect 154166 79834 154218 79840
rect 154270 79778 154298 80036
rect 153994 79750 154068 79778
rect 153936 79688 153988 79694
rect 153936 79630 153988 79636
rect 153948 76673 153976 79630
rect 154040 78577 154068 79750
rect 154120 79756 154172 79762
rect 154120 79698 154172 79704
rect 154224 79750 154298 79778
rect 154362 79778 154390 80036
rect 154454 79937 154482 80036
rect 154546 79966 154574 80036
rect 154638 79966 154666 80036
rect 154730 79966 154758 80036
rect 154534 79960 154586 79966
rect 154440 79928 154496 79937
rect 154534 79902 154586 79908
rect 154626 79960 154678 79966
rect 154626 79902 154678 79908
rect 154718 79960 154770 79966
rect 154718 79902 154770 79908
rect 154440 79863 154496 79872
rect 154822 79812 154850 80036
rect 154578 79792 154634 79801
rect 154362 79750 154436 79778
rect 154132 78674 154160 79698
rect 154224 79665 154252 79750
rect 154304 79688 154356 79694
rect 154210 79656 154266 79665
rect 154304 79630 154356 79636
rect 154210 79591 154266 79600
rect 154316 79529 154344 79630
rect 154302 79520 154358 79529
rect 154302 79455 154358 79464
rect 154210 79384 154266 79393
rect 154210 79319 154266 79328
rect 154120 78668 154172 78674
rect 154120 78610 154172 78616
rect 154026 78568 154082 78577
rect 154026 78503 154082 78512
rect 154118 77888 154174 77897
rect 154118 77823 154174 77832
rect 153934 76664 153990 76673
rect 153934 76599 153990 76608
rect 153936 76424 153988 76430
rect 153936 76366 153988 76372
rect 153948 75614 153976 76366
rect 153936 75608 153988 75614
rect 153936 75550 153988 75556
rect 153844 75268 153896 75274
rect 153844 75210 153896 75216
rect 154132 75154 154160 77823
rect 153764 75126 154160 75154
rect 153660 70236 153712 70242
rect 153660 70178 153712 70184
rect 153568 70032 153620 70038
rect 153568 69974 153620 69980
rect 153108 60036 153160 60042
rect 153108 59978 153160 59984
rect 153764 20194 153792 75126
rect 154120 75064 154172 75070
rect 154120 75006 154172 75012
rect 154028 74520 154080 74526
rect 154028 74462 154080 74468
rect 153844 70372 153896 70378
rect 153844 70314 153896 70320
rect 153752 20188 153804 20194
rect 153752 20130 153804 20136
rect 153016 16176 153068 16182
rect 153016 16118 153068 16124
rect 153856 13394 153884 70314
rect 153936 70032 153988 70038
rect 153936 69974 153988 69980
rect 153948 14754 153976 69974
rect 154040 25838 154068 74462
rect 154132 70174 154160 75006
rect 154224 70394 154252 79319
rect 154304 75744 154356 75750
rect 154304 75686 154356 75692
rect 154316 75002 154344 75686
rect 154408 75070 154436 79750
rect 154776 79784 154850 79812
rect 154578 79727 154634 79736
rect 154672 79756 154724 79762
rect 154488 79688 154540 79694
rect 154488 79630 154540 79636
rect 154500 78577 154528 79630
rect 154486 78568 154542 78577
rect 154486 78503 154542 78512
rect 154488 78464 154540 78470
rect 154592 78452 154620 79727
rect 154672 79698 154724 79704
rect 154684 78554 154712 79698
rect 154776 79354 154804 79784
rect 154914 79744 154942 80036
rect 155006 79937 155034 80036
rect 154992 79928 155048 79937
rect 154992 79863 155048 79872
rect 155098 79812 155126 80036
rect 155190 79966 155218 80036
rect 155282 79966 155310 80036
rect 155178 79960 155230 79966
rect 155178 79902 155230 79908
rect 155270 79960 155322 79966
rect 155270 79902 155322 79908
rect 155270 79824 155322 79830
rect 155098 79784 155172 79812
rect 154868 79716 154942 79744
rect 154764 79348 154816 79354
rect 154764 79290 154816 79296
rect 154684 78526 154804 78554
rect 154592 78424 154712 78452
rect 154488 78406 154540 78412
rect 154396 75064 154448 75070
rect 154396 75006 154448 75012
rect 154304 74996 154356 75002
rect 154304 74938 154356 74944
rect 154500 70394 154528 78406
rect 154578 76936 154634 76945
rect 154578 76871 154634 76880
rect 154224 70366 154344 70394
rect 154212 70236 154264 70242
rect 154212 70178 154264 70184
rect 154120 70168 154172 70174
rect 154120 70110 154172 70116
rect 154028 25832 154080 25838
rect 154028 25774 154080 25780
rect 154132 24342 154160 70110
rect 154224 32638 154252 70178
rect 154316 46374 154344 70366
rect 154408 70366 154528 70394
rect 154304 46368 154356 46374
rect 154304 46310 154356 46316
rect 154212 32632 154264 32638
rect 154212 32574 154264 32580
rect 154120 24336 154172 24342
rect 154120 24278 154172 24284
rect 154408 20262 154436 70366
rect 154592 68241 154620 76871
rect 154578 68232 154634 68241
rect 154578 68167 154634 68176
rect 154684 38214 154712 78424
rect 154776 70394 154804 78526
rect 154868 77382 154896 79716
rect 155040 79688 155092 79694
rect 155040 79630 155092 79636
rect 154856 77376 154908 77382
rect 154856 77318 154908 77324
rect 155052 73778 155080 79630
rect 155144 78577 155172 79784
rect 155222 79792 155270 79801
rect 155278 79766 155322 79772
rect 155278 79750 155310 79766
rect 155222 79727 155278 79736
rect 155224 79688 155276 79694
rect 155374 79676 155402 80036
rect 155466 79812 155494 80036
rect 155558 79937 155586 80036
rect 155544 79928 155600 79937
rect 155544 79863 155600 79872
rect 155650 79830 155678 80036
rect 155742 79966 155770 80036
rect 155730 79960 155782 79966
rect 155834 79937 155862 80036
rect 155926 79966 155954 80036
rect 155914 79960 155966 79966
rect 155730 79902 155782 79908
rect 155820 79928 155876 79937
rect 155914 79902 155966 79908
rect 155820 79863 155876 79872
rect 155638 79824 155690 79830
rect 155466 79784 155540 79812
rect 155374 79648 155448 79676
rect 155224 79630 155276 79636
rect 155130 78568 155186 78577
rect 155130 78503 155186 78512
rect 155236 74746 155264 79630
rect 155316 79484 155368 79490
rect 155316 79426 155368 79432
rect 155328 75041 155356 79426
rect 155420 77897 155448 79648
rect 155406 77888 155462 77897
rect 155406 77823 155462 77832
rect 155512 76974 155540 79784
rect 155834 79812 155862 79863
rect 156018 79812 156046 80036
rect 156110 79966 156138 80036
rect 156098 79960 156150 79966
rect 156098 79902 156150 79908
rect 155834 79784 155908 79812
rect 156018 79784 156092 79812
rect 155638 79766 155690 79772
rect 155590 79656 155646 79665
rect 155590 79591 155646 79600
rect 155684 79620 155736 79626
rect 155500 76968 155552 76974
rect 155500 76910 155552 76916
rect 155314 75032 155370 75041
rect 155370 74990 155448 75018
rect 155314 74967 155370 74976
rect 155236 74718 155356 74746
rect 155328 73817 155356 74718
rect 155314 73808 155370 73817
rect 155040 73772 155092 73778
rect 155314 73743 155370 73752
rect 155040 73714 155092 73720
rect 154776 70366 155264 70394
rect 155236 70310 155264 70366
rect 155224 70304 155276 70310
rect 155224 70246 155276 70252
rect 155236 49094 155264 70246
rect 155328 60110 155356 73743
rect 155316 60104 155368 60110
rect 155316 60046 155368 60052
rect 155224 49088 155276 49094
rect 155224 49030 155276 49036
rect 155420 42362 155448 74990
rect 155604 74050 155632 79591
rect 155684 79562 155736 79568
rect 155696 74225 155724 79562
rect 155774 79520 155830 79529
rect 155774 79455 155830 79464
rect 155682 74216 155738 74225
rect 155682 74151 155738 74160
rect 155592 74044 155644 74050
rect 155592 73986 155644 73992
rect 155696 73930 155724 74151
rect 155512 73902 155724 73930
rect 155408 42356 155460 42362
rect 155408 42298 155460 42304
rect 154672 38208 154724 38214
rect 154672 38150 154724 38156
rect 154580 37936 154632 37942
rect 154580 37878 154632 37884
rect 154396 20256 154448 20262
rect 154396 20198 154448 20204
rect 154592 16574 154620 37878
rect 155512 36718 155540 73902
rect 155684 73772 155736 73778
rect 155684 73714 155736 73720
rect 155696 73030 155724 73714
rect 155684 73024 155736 73030
rect 155684 72966 155736 72972
rect 155500 36712 155552 36718
rect 155500 36654 155552 36660
rect 155696 19990 155724 72966
rect 155788 20126 155816 79455
rect 155776 20120 155828 20126
rect 155776 20062 155828 20068
rect 155684 19984 155736 19990
rect 155684 19926 155736 19932
rect 155880 18834 155908 79784
rect 156064 79506 156092 79784
rect 156202 79744 156230 80036
rect 156294 79966 156322 80036
rect 156282 79960 156334 79966
rect 156282 79902 156334 79908
rect 156282 79824 156334 79830
rect 156386 79801 156414 80036
rect 156478 79966 156506 80036
rect 156570 79966 156598 80036
rect 156466 79960 156518 79966
rect 156466 79902 156518 79908
rect 156558 79960 156610 79966
rect 156558 79902 156610 79908
rect 156662 79801 156690 80036
rect 156282 79766 156334 79772
rect 156372 79792 156428 79801
rect 155972 79478 156092 79506
rect 156156 79716 156230 79744
rect 155972 73001 156000 79478
rect 156052 79416 156104 79422
rect 156052 79358 156104 79364
rect 155958 72992 156014 73001
rect 155958 72927 156014 72936
rect 155960 72888 156012 72894
rect 155960 72830 156012 72836
rect 155972 51814 156000 72830
rect 156064 70281 156092 79358
rect 156156 77654 156184 79716
rect 156294 79676 156322 79766
rect 156648 79792 156704 79801
rect 156372 79727 156428 79736
rect 156616 79736 156648 79744
rect 156616 79727 156704 79736
rect 156754 79744 156782 80036
rect 156846 79966 156874 80036
rect 156938 79966 156966 80036
rect 156834 79960 156886 79966
rect 156834 79902 156886 79908
rect 156926 79960 156978 79966
rect 157030 79937 157058 80036
rect 156926 79902 156978 79908
rect 157016 79928 157072 79937
rect 157016 79863 157072 79872
rect 156972 79824 157024 79830
rect 156972 79766 157024 79772
rect 156248 79648 156322 79676
rect 156616 79716 156690 79727
rect 156754 79716 156828 79744
rect 156248 77874 156276 79648
rect 156512 79620 156564 79626
rect 156512 79562 156564 79568
rect 156328 79552 156380 79558
rect 156328 79494 156380 79500
rect 156340 78169 156368 79494
rect 156420 79484 156472 79490
rect 156420 79426 156472 79432
rect 156326 78160 156382 78169
rect 156326 78095 156382 78104
rect 156432 77994 156460 79426
rect 156420 77988 156472 77994
rect 156420 77930 156472 77936
rect 156524 77897 156552 79562
rect 156510 77888 156566 77897
rect 156248 77846 156460 77874
rect 156144 77648 156196 77654
rect 156144 77590 156196 77596
rect 156326 77616 156382 77625
rect 156326 77551 156382 77560
rect 156340 73137 156368 77551
rect 156326 73128 156382 73137
rect 156326 73063 156382 73072
rect 156050 70272 156106 70281
rect 156050 70207 156106 70216
rect 156064 69873 156092 70207
rect 156050 69864 156106 69873
rect 156050 69799 156106 69808
rect 155960 51808 156012 51814
rect 155960 51750 156012 51756
rect 156340 43586 156368 73063
rect 156432 71738 156460 77846
rect 156510 77823 156566 77832
rect 156616 72826 156644 79716
rect 156696 79620 156748 79626
rect 156696 79562 156748 79568
rect 156708 77178 156736 79562
rect 156800 78441 156828 79716
rect 156984 79665 157012 79766
rect 157122 79676 157150 80036
rect 157214 79937 157242 80036
rect 157306 79966 157334 80036
rect 157294 79960 157346 79966
rect 157200 79928 157256 79937
rect 157294 79902 157346 79908
rect 157200 79863 157256 79872
rect 157214 79812 157242 79863
rect 157398 79812 157426 80036
rect 157214 79784 157288 79812
rect 156970 79656 157026 79665
rect 156892 79614 156970 79642
rect 156786 78432 156842 78441
rect 156786 78367 156842 78376
rect 156892 78316 156920 79614
rect 156970 79591 157026 79600
rect 157076 79648 157150 79676
rect 156972 79552 157024 79558
rect 156972 79494 157024 79500
rect 156984 78713 157012 79494
rect 156970 78704 157026 78713
rect 156970 78639 157026 78648
rect 156800 78288 156920 78316
rect 156696 77172 156748 77178
rect 156696 77114 156748 77120
rect 156604 72820 156656 72826
rect 156604 72762 156656 72768
rect 156800 72706 156828 78288
rect 156880 77172 156932 77178
rect 156880 77114 156932 77120
rect 156524 72678 156828 72706
rect 156420 71732 156472 71738
rect 156420 71674 156472 71680
rect 156524 70394 156552 72678
rect 156602 72312 156658 72321
rect 156602 72247 156658 72256
rect 156432 70366 156552 70394
rect 156328 43580 156380 43586
rect 156328 43522 156380 43528
rect 155868 18828 155920 18834
rect 155868 18770 155920 18776
rect 154592 16546 155448 16574
rect 153936 14748 153988 14754
rect 153936 14690 153988 14696
rect 153844 13388 153896 13394
rect 153844 13330 153896 13336
rect 152464 10600 152516 10606
rect 152464 10542 152516 10548
rect 152096 5024 152148 5030
rect 152096 4966 152148 4972
rect 153016 4072 153068 4078
rect 153016 4014 153068 4020
rect 151832 3454 151952 3482
rect 151832 480 151860 3454
rect 153028 480 153056 4014
rect 154212 3188 154264 3194
rect 154212 3130 154264 3136
rect 154224 480 154252 3130
rect 155420 480 155448 16546
rect 156432 6458 156460 70366
rect 156616 6914 156644 72247
rect 156892 71777 156920 77114
rect 156984 72894 157012 78639
rect 157076 76809 157104 79648
rect 157062 76800 157118 76809
rect 157062 76735 157118 76744
rect 156972 72888 157024 72894
rect 156972 72830 157024 72836
rect 156878 71768 156934 71777
rect 156696 71732 156748 71738
rect 156878 71703 156934 71712
rect 156696 71674 156748 71680
rect 156708 10538 156736 71674
rect 156786 69864 156842 69873
rect 156786 69799 156842 69808
rect 156800 14686 156828 69799
rect 156892 35494 156920 71703
rect 157076 40934 157104 76735
rect 157154 72992 157210 73001
rect 157154 72927 157210 72936
rect 157064 40928 157116 40934
rect 157064 40870 157116 40876
rect 156880 35488 156932 35494
rect 156880 35430 156932 35436
rect 157168 31346 157196 72927
rect 157260 72758 157288 79784
rect 157352 79784 157426 79812
rect 157352 73166 157380 79784
rect 157490 79744 157518 80036
rect 157582 79830 157610 80036
rect 157674 79966 157702 80036
rect 157662 79960 157714 79966
rect 157766 79937 157794 80036
rect 157662 79902 157714 79908
rect 157752 79928 157808 79937
rect 157752 79863 157808 79872
rect 157570 79824 157622 79830
rect 157858 79812 157886 80036
rect 157570 79766 157622 79772
rect 157706 79792 157762 79801
rect 157444 79716 157518 79744
rect 157706 79727 157762 79736
rect 157812 79784 157886 79812
rect 157444 77858 157472 79716
rect 157616 79552 157668 79558
rect 157616 79494 157668 79500
rect 157524 79484 157576 79490
rect 157524 79426 157576 79432
rect 157432 77852 157484 77858
rect 157432 77794 157484 77800
rect 157444 77761 157472 77794
rect 157430 77752 157486 77761
rect 157430 77687 157486 77696
rect 157430 75304 157486 75313
rect 157430 75239 157486 75248
rect 157340 73160 157392 73166
rect 157340 73102 157392 73108
rect 157248 72752 157300 72758
rect 157248 72694 157300 72700
rect 157444 72457 157472 75239
rect 157536 73098 157564 79426
rect 157628 79082 157656 79494
rect 157616 79076 157668 79082
rect 157616 79018 157668 79024
rect 157616 78940 157668 78946
rect 157616 78882 157668 78888
rect 157524 73092 157576 73098
rect 157524 73034 157576 73040
rect 157628 72622 157656 78882
rect 157720 72690 157748 79727
rect 157812 79665 157840 79784
rect 157950 79744 157978 80036
rect 158042 79830 158070 80036
rect 158030 79824 158082 79830
rect 158030 79766 158082 79772
rect 158134 79778 158162 80036
rect 158226 79898 158254 80036
rect 158318 79966 158346 80036
rect 158306 79960 158358 79966
rect 158306 79902 158358 79908
rect 158214 79892 158266 79898
rect 158214 79834 158266 79840
rect 158410 79812 158438 80036
rect 158502 79898 158530 80036
rect 158594 79937 158622 80036
rect 158580 79928 158636 79937
rect 158490 79892 158542 79898
rect 158686 79898 158714 80036
rect 158778 79898 158806 80036
rect 158580 79863 158636 79872
rect 158674 79892 158726 79898
rect 158490 79834 158542 79840
rect 158364 79784 158438 79812
rect 158364 79778 158392 79784
rect 158134 79750 158208 79778
rect 157904 79716 157978 79744
rect 157798 79656 157854 79665
rect 157798 79591 157854 79600
rect 157798 79520 157854 79529
rect 157798 79455 157800 79464
rect 157852 79455 157854 79464
rect 157800 79426 157852 79432
rect 157812 78946 157840 79426
rect 157800 78940 157852 78946
rect 157800 78882 157852 78888
rect 157800 77852 157852 77858
rect 157800 77794 157852 77800
rect 157708 72684 157760 72690
rect 157708 72626 157760 72632
rect 157616 72616 157668 72622
rect 157616 72558 157668 72564
rect 157430 72448 157486 72457
rect 157430 72383 157486 72392
rect 157156 31340 157208 31346
rect 157156 31282 157208 31288
rect 157812 21622 157840 77794
rect 157904 77294 157932 79716
rect 158076 79688 158128 79694
rect 158074 79656 158076 79665
rect 158128 79656 158130 79665
rect 158074 79591 158130 79600
rect 157904 77266 158024 77294
rect 157996 74474 158024 77266
rect 158088 77194 158116 79591
rect 158180 78713 158208 79750
rect 158272 79750 158392 79778
rect 158166 78704 158222 78713
rect 158166 78639 158222 78648
rect 158088 77166 158208 77194
rect 157996 74446 158116 74474
rect 157982 74352 158038 74361
rect 157982 74287 158038 74296
rect 157996 53174 158024 74287
rect 158088 74089 158116 74446
rect 158180 74202 158208 77166
rect 158272 74361 158300 79750
rect 158594 79744 158622 79863
rect 158674 79834 158726 79840
rect 158766 79892 158818 79898
rect 158766 79834 158818 79840
rect 158870 79801 158898 80036
rect 158456 79716 158622 79744
rect 158856 79792 158912 79801
rect 158856 79727 158912 79736
rect 158962 79744 158990 80036
rect 159054 79966 159082 80036
rect 159146 79966 159174 80036
rect 159042 79960 159094 79966
rect 159042 79902 159094 79908
rect 159134 79960 159186 79966
rect 159134 79902 159186 79908
rect 159238 79744 159266 80036
rect 158352 79688 158404 79694
rect 158352 79630 158404 79636
rect 158364 77450 158392 79630
rect 158352 77444 158404 77450
rect 158352 77386 158404 77392
rect 158258 74352 158314 74361
rect 158258 74287 158314 74296
rect 158180 74174 158392 74202
rect 158074 74080 158130 74089
rect 158074 74015 158130 74024
rect 158260 73160 158312 73166
rect 158260 73102 158312 73108
rect 158272 72486 158300 73102
rect 158260 72480 158312 72486
rect 158260 72422 158312 72428
rect 157984 53168 158036 53174
rect 157984 53110 158036 53116
rect 158272 29918 158300 72422
rect 158260 29912 158312 29918
rect 158260 29854 158312 29860
rect 157800 21616 157852 21622
rect 157800 21558 157852 21564
rect 158364 21554 158392 74174
rect 158352 21548 158404 21554
rect 158352 21490 158404 21496
rect 158456 21486 158484 79716
rect 158870 79676 158898 79727
rect 158962 79716 159036 79744
rect 158824 79648 158898 79676
rect 158536 79620 158588 79626
rect 158536 79562 158588 79568
rect 158628 79620 158680 79626
rect 158628 79562 158680 79568
rect 158548 78713 158576 79562
rect 158534 78704 158590 78713
rect 158534 78639 158590 78648
rect 158640 77897 158668 79562
rect 158718 79248 158774 79257
rect 158718 79183 158774 79192
rect 158626 77888 158682 77897
rect 158626 77823 158682 77832
rect 158628 77376 158680 77382
rect 158628 77318 158680 77324
rect 158640 76022 158668 77318
rect 158628 76016 158680 76022
rect 158628 75958 158680 75964
rect 158626 74080 158682 74089
rect 158626 74015 158682 74024
rect 158640 73817 158668 74015
rect 158626 73808 158682 73817
rect 158626 73743 158682 73752
rect 158536 73092 158588 73098
rect 158536 73034 158588 73040
rect 158548 72418 158576 73034
rect 158536 72412 158588 72418
rect 158536 72354 158588 72360
rect 158444 21480 158496 21486
rect 158444 21422 158496 21428
rect 156788 14680 156840 14686
rect 156788 14622 156840 14628
rect 158548 13326 158576 72354
rect 158536 13320 158588 13326
rect 158536 13262 158588 13268
rect 156696 10532 156748 10538
rect 156696 10474 156748 10480
rect 158640 9246 158668 73743
rect 158732 21418 158760 79183
rect 158824 78470 158852 79648
rect 158904 79552 158956 79558
rect 158904 79494 158956 79500
rect 158812 78464 158864 78470
rect 158812 78406 158864 78412
rect 158916 75426 158944 79494
rect 158824 75398 158944 75426
rect 158824 71670 158852 75398
rect 158904 75268 158956 75274
rect 158904 75210 158956 75216
rect 158812 71664 158864 71670
rect 158812 71606 158864 71612
rect 158812 71528 158864 71534
rect 158812 71470 158864 71476
rect 158824 38146 158852 71470
rect 158916 60722 158944 75210
rect 159008 63510 159036 79716
rect 159192 79716 159266 79744
rect 159088 79484 159140 79490
rect 159088 79426 159140 79432
rect 159100 79257 159128 79426
rect 159086 79248 159142 79257
rect 159086 79183 159142 79192
rect 159192 75274 159220 79716
rect 159330 79608 159358 80036
rect 159422 79801 159450 80036
rect 159514 79971 159542 80036
rect 159500 79962 159556 79971
rect 159606 79966 159634 80036
rect 159500 79897 159556 79906
rect 159594 79960 159646 79966
rect 159698 79937 159726 80036
rect 159594 79902 159646 79908
rect 159684 79928 159740 79937
rect 159790 79898 159818 80036
rect 159684 79863 159740 79872
rect 159778 79892 159830 79898
rect 159778 79834 159830 79840
rect 159548 79824 159600 79830
rect 159408 79792 159464 79801
rect 159548 79766 159600 79772
rect 159464 79736 159496 79744
rect 159408 79727 159496 79736
rect 159422 79716 159496 79727
rect 159284 79580 159358 79608
rect 159180 75268 159232 75274
rect 159180 75210 159232 75216
rect 159284 70394 159312 79580
rect 159364 79484 159416 79490
rect 159364 79426 159416 79432
rect 159376 77790 159404 79426
rect 159364 77784 159416 77790
rect 159364 77726 159416 77732
rect 159376 71534 159404 77726
rect 159468 77246 159496 79716
rect 159456 77240 159508 77246
rect 159456 77182 159508 77188
rect 159560 75914 159588 79766
rect 159882 79744 159910 80036
rect 159974 79971 160002 80036
rect 159960 79962 160016 79971
rect 159960 79897 160016 79906
rect 160066 79744 160094 80036
rect 159836 79716 159910 79744
rect 160020 79716 160094 79744
rect 159638 79656 159694 79665
rect 159638 79591 159694 79600
rect 159652 79558 159680 79591
rect 159640 79552 159692 79558
rect 159640 79494 159692 79500
rect 159732 79416 159784 79422
rect 159732 79358 159784 79364
rect 159560 75886 159680 75914
rect 159652 71738 159680 75886
rect 159744 74066 159772 79358
rect 159836 77110 159864 79716
rect 159916 79552 159968 79558
rect 159916 79494 159968 79500
rect 159824 77104 159876 77110
rect 159824 77046 159876 77052
rect 159744 74038 159864 74066
rect 159836 71777 159864 74038
rect 159822 71768 159878 71777
rect 159640 71732 159692 71738
rect 159822 71703 159878 71712
rect 159640 71674 159692 71680
rect 159732 71664 159784 71670
rect 159732 71606 159784 71612
rect 159364 71528 159416 71534
rect 159364 71470 159416 71476
rect 159744 71262 159772 71606
rect 159732 71256 159784 71262
rect 159732 71198 159784 71204
rect 159100 70366 159312 70394
rect 159100 66230 159128 70366
rect 159088 66224 159140 66230
rect 159088 66166 159140 66172
rect 158996 63504 159048 63510
rect 158996 63446 159048 63452
rect 158904 60716 158956 60722
rect 158904 60658 158956 60664
rect 158812 38140 158864 38146
rect 158812 38082 158864 38088
rect 159744 35426 159772 71198
rect 159732 35420 159784 35426
rect 159732 35362 159784 35368
rect 159836 28490 159864 71703
rect 159824 28484 159876 28490
rect 159824 28426 159876 28432
rect 159928 22982 159956 79494
rect 160020 78441 160048 79716
rect 160158 79642 160186 80036
rect 160250 79801 160278 80036
rect 160342 79937 160370 80036
rect 160434 79966 160462 80036
rect 160526 79966 160554 80036
rect 160422 79960 160474 79966
rect 160328 79928 160384 79937
rect 160422 79902 160474 79908
rect 160514 79960 160566 79966
rect 160514 79902 160566 79908
rect 160328 79863 160384 79872
rect 160376 79824 160428 79830
rect 160236 79792 160292 79801
rect 160376 79766 160428 79772
rect 160236 79727 160292 79736
rect 160158 79614 160324 79642
rect 160190 79112 160246 79121
rect 160190 79047 160246 79056
rect 160006 78432 160062 78441
rect 160006 78367 160062 78376
rect 160008 71732 160060 71738
rect 160008 71674 160060 71680
rect 160020 70990 160048 71674
rect 160008 70984 160060 70990
rect 160008 70926 160060 70932
rect 159916 22976 159968 22982
rect 159916 22918 159968 22924
rect 158720 21412 158772 21418
rect 158720 21354 158772 21360
rect 158718 21312 158774 21321
rect 158718 21247 158774 21256
rect 158732 16574 158760 21247
rect 158732 16546 158944 16574
rect 158628 9240 158680 9246
rect 158628 9182 158680 9188
rect 156616 6886 156736 6914
rect 156420 6452 156472 6458
rect 156420 6394 156472 6400
rect 156708 3942 156736 6886
rect 157800 4004 157852 4010
rect 157800 3946 157852 3952
rect 156604 3936 156656 3942
rect 156604 3878 156656 3884
rect 156696 3936 156748 3942
rect 156696 3878 156748 3884
rect 156616 480 156644 3878
rect 157812 480 157840 3946
rect 158916 480 158944 16546
rect 160020 7750 160048 70926
rect 160100 70916 160152 70922
rect 160100 70858 160152 70864
rect 160112 16046 160140 70858
rect 160204 62830 160232 79047
rect 160296 71670 160324 79614
rect 160388 73166 160416 79766
rect 160468 79756 160520 79762
rect 160618 79744 160646 80036
rect 160710 79898 160738 80036
rect 160802 79898 160830 80036
rect 160894 79966 160922 80036
rect 160882 79960 160934 79966
rect 160882 79902 160934 79908
rect 160698 79892 160750 79898
rect 160698 79834 160750 79840
rect 160790 79892 160842 79898
rect 160790 79834 160842 79840
rect 160468 79698 160520 79704
rect 160572 79716 160646 79744
rect 160742 79792 160798 79801
rect 160742 79727 160744 79736
rect 160480 78826 160508 79698
rect 160572 79121 160600 79716
rect 160796 79727 160798 79736
rect 160986 79744 161014 80036
rect 161078 79966 161106 80036
rect 161170 79966 161198 80036
rect 161262 79966 161290 80036
rect 161066 79960 161118 79966
rect 161066 79902 161118 79908
rect 161158 79960 161210 79966
rect 161158 79902 161210 79908
rect 161250 79960 161302 79966
rect 161250 79902 161302 79908
rect 161354 79830 161382 80036
rect 161446 79937 161474 80036
rect 161432 79928 161488 79937
rect 161432 79863 161488 79872
rect 161342 79824 161394 79830
rect 161202 79792 161258 79801
rect 161112 79756 161164 79762
rect 160986 79716 161060 79744
rect 160744 79698 160796 79704
rect 160652 79620 160704 79626
rect 160652 79562 160704 79568
rect 160664 79150 160692 79562
rect 160652 79144 160704 79150
rect 160558 79112 160614 79121
rect 160652 79086 160704 79092
rect 160558 79047 160614 79056
rect 160480 78798 160600 78826
rect 160466 78704 160522 78713
rect 160466 78639 160522 78648
rect 160376 73160 160428 73166
rect 160376 73102 160428 73108
rect 160284 71664 160336 71670
rect 160284 71606 160336 71612
rect 160480 71058 160508 78639
rect 160572 78033 160600 78798
rect 160558 78024 160614 78033
rect 160558 77959 160614 77968
rect 160468 71052 160520 71058
rect 160468 70994 160520 71000
rect 160572 70394 160600 77959
rect 160664 75914 160692 79086
rect 160756 77382 160784 79698
rect 160836 79688 160888 79694
rect 160836 79630 160888 79636
rect 160926 79656 160982 79665
rect 160744 77376 160796 77382
rect 160848 77353 160876 79630
rect 160926 79591 160928 79600
rect 160980 79591 160982 79600
rect 160928 79562 160980 79568
rect 160940 78266 160968 79562
rect 160928 78260 160980 78266
rect 160928 78202 160980 78208
rect 160744 77318 160796 77324
rect 160834 77344 160890 77353
rect 160834 77279 160890 77288
rect 161032 77178 161060 79716
rect 161342 79766 161394 79772
rect 161202 79727 161258 79736
rect 161112 79698 161164 79704
rect 161124 77353 161152 79698
rect 161216 79694 161244 79727
rect 161204 79688 161256 79694
rect 161538 79676 161566 80036
rect 161630 79966 161658 80036
rect 161618 79960 161670 79966
rect 161722 79937 161750 80036
rect 161618 79902 161670 79908
rect 161708 79928 161764 79937
rect 161708 79863 161764 79872
rect 161664 79824 161716 79830
rect 161814 79778 161842 80036
rect 161906 79830 161934 80036
rect 161998 79966 162026 80036
rect 161986 79960 162038 79966
rect 161986 79902 162038 79908
rect 161664 79766 161716 79772
rect 161204 79630 161256 79636
rect 161492 79648 161566 79676
rect 161110 77344 161166 77353
rect 161110 77279 161166 77288
rect 161020 77172 161072 77178
rect 161020 77114 161072 77120
rect 160836 76424 160888 76430
rect 160836 76366 160888 76372
rect 160664 75886 160784 75914
rect 160756 70922 160784 75886
rect 160848 71738 160876 76366
rect 161112 73160 161164 73166
rect 161112 73102 161164 73108
rect 161124 72282 161152 73102
rect 161112 72276 161164 72282
rect 161112 72218 161164 72224
rect 160836 71732 160888 71738
rect 160836 71674 160888 71680
rect 161020 71664 161072 71670
rect 161020 71606 161072 71612
rect 160744 70916 160796 70922
rect 160744 70858 160796 70864
rect 160572 70366 160784 70394
rect 160192 62824 160244 62830
rect 160192 62766 160244 62772
rect 160756 39574 160784 70366
rect 160744 39568 160796 39574
rect 160744 39510 160796 39516
rect 161032 32570 161060 71606
rect 161020 32564 161072 32570
rect 161020 32506 161072 32512
rect 161124 16114 161152 72218
rect 161216 20058 161244 79630
rect 161296 79620 161348 79626
rect 161296 79562 161348 79568
rect 161308 76430 161336 79562
rect 161492 78198 161520 79648
rect 161572 79416 161624 79422
rect 161572 79358 161624 79364
rect 161480 78192 161532 78198
rect 161480 78134 161532 78140
rect 161480 77988 161532 77994
rect 161480 77930 161532 77936
rect 161388 77376 161440 77382
rect 161388 77318 161440 77324
rect 161296 76424 161348 76430
rect 161296 76366 161348 76372
rect 161296 71732 161348 71738
rect 161296 71674 161348 71680
rect 161308 71398 161336 71674
rect 161296 71392 161348 71398
rect 161296 71334 161348 71340
rect 161204 20052 161256 20058
rect 161204 19994 161256 20000
rect 161112 16108 161164 16114
rect 161112 16050 161164 16056
rect 160100 16040 160152 16046
rect 160100 15982 160152 15988
rect 160098 15872 160154 15881
rect 160098 15807 160154 15816
rect 160008 7744 160060 7750
rect 160008 7686 160060 7692
rect 160112 480 160140 15807
rect 161308 6390 161336 71334
rect 161400 9178 161428 77318
rect 161492 68950 161520 77930
rect 161480 68944 161532 68950
rect 161480 68886 161532 68892
rect 161584 45014 161612 79358
rect 161676 78849 161704 79766
rect 161768 79750 161842 79778
rect 161894 79824 161946 79830
rect 161894 79766 161946 79772
rect 161662 78840 161718 78849
rect 161662 78775 161718 78784
rect 161676 77382 161704 78775
rect 161664 77376 161716 77382
rect 161664 77318 161716 77324
rect 161664 77240 161716 77246
rect 161664 77182 161716 77188
rect 161676 73982 161704 77182
rect 161768 76702 161796 79750
rect 162090 79744 162118 80036
rect 162182 79966 162210 80036
rect 162170 79960 162222 79966
rect 162170 79902 162222 79908
rect 162274 79778 162302 80036
rect 162366 79898 162394 80036
rect 162458 79937 162486 80036
rect 162444 79928 162500 79937
rect 162354 79892 162406 79898
rect 162550 79898 162578 80036
rect 162642 79898 162670 80036
rect 162734 79937 162762 80036
rect 162720 79928 162776 79937
rect 162444 79863 162500 79872
rect 162538 79892 162590 79898
rect 162354 79834 162406 79840
rect 162538 79834 162590 79840
rect 162630 79892 162682 79898
rect 162826 79898 162854 80036
rect 162918 79971 162946 80036
rect 162904 79962 162960 79971
rect 163010 79966 163038 80036
rect 163102 79966 163130 80036
rect 162720 79863 162776 79872
rect 162814 79892 162866 79898
rect 162904 79897 162960 79906
rect 162998 79960 163050 79966
rect 162998 79902 163050 79908
rect 163090 79960 163142 79966
rect 163090 79902 163142 79908
rect 162630 79834 162682 79840
rect 162814 79834 162866 79840
rect 163194 79830 163222 80036
rect 163286 79898 163314 80036
rect 163378 79966 163406 80036
rect 163366 79960 163418 79966
rect 163366 79902 163418 79908
rect 163274 79892 163326 79898
rect 163274 79834 163326 79840
rect 163470 79830 163498 80036
rect 163182 79824 163234 79830
rect 162858 79792 162914 79801
rect 162274 79750 162348 79778
rect 162090 79716 162164 79744
rect 161848 79688 161900 79694
rect 161848 79630 161900 79636
rect 161860 79121 161888 79630
rect 161940 79620 161992 79626
rect 161940 79562 161992 79568
rect 161846 79112 161902 79121
rect 161846 79047 161902 79056
rect 161846 78976 161902 78985
rect 161952 78928 161980 79562
rect 161902 78920 161980 78928
rect 161846 78911 161980 78920
rect 161860 78900 161980 78911
rect 161756 76696 161808 76702
rect 161756 76638 161808 76644
rect 161756 76492 161808 76498
rect 161756 76434 161808 76440
rect 161664 73976 161716 73982
rect 161664 73918 161716 73924
rect 161768 70394 161796 76434
rect 161676 70366 161796 70394
rect 161860 70394 161888 78900
rect 162032 78192 162084 78198
rect 162032 78134 162084 78140
rect 161940 76696 161992 76702
rect 161940 76638 161992 76644
rect 161952 71738 161980 76638
rect 162044 73154 162072 78134
rect 162136 74746 162164 79716
rect 162216 79688 162268 79694
rect 162216 79630 162268 79636
rect 162228 79529 162256 79630
rect 162214 79520 162270 79529
rect 162214 79455 162270 79464
rect 162228 78849 162256 79455
rect 162214 78840 162270 78849
rect 162214 78775 162270 78784
rect 162216 77648 162268 77654
rect 162216 77590 162268 77596
rect 162228 77314 162256 77590
rect 162216 77308 162268 77314
rect 162216 77250 162268 77256
rect 162320 76537 162348 79750
rect 162584 79756 162636 79762
rect 162584 79698 162636 79704
rect 162676 79756 162728 79762
rect 163182 79766 163234 79772
rect 163458 79824 163510 79830
rect 163458 79766 163510 79772
rect 162858 79727 162914 79736
rect 162952 79756 163004 79762
rect 162676 79698 162728 79704
rect 162490 79656 162546 79665
rect 162400 79620 162452 79626
rect 162490 79591 162546 79600
rect 162400 79562 162452 79568
rect 162306 76528 162362 76537
rect 162412 76498 162440 79562
rect 162306 76463 162362 76472
rect 162400 76492 162452 76498
rect 162400 76434 162452 76440
rect 162504 75018 162532 79591
rect 162596 75993 162624 79698
rect 162688 79529 162716 79698
rect 162766 79656 162822 79665
rect 162766 79591 162822 79600
rect 162674 79520 162730 79529
rect 162674 79455 162730 79464
rect 162582 75984 162638 75993
rect 162582 75919 162638 75928
rect 162688 75138 162716 79455
rect 162676 75132 162728 75138
rect 162676 75074 162728 75080
rect 162504 74990 162716 75018
rect 162136 74718 162440 74746
rect 162044 73126 162164 73154
rect 161940 71732 161992 71738
rect 161940 71674 161992 71680
rect 162136 71466 162164 73126
rect 162124 71460 162176 71466
rect 162124 71402 162176 71408
rect 162136 70394 162164 71402
rect 162412 71330 162440 74718
rect 162584 71732 162636 71738
rect 162584 71674 162636 71680
rect 162596 71602 162624 71674
rect 162584 71596 162636 71602
rect 162584 71538 162636 71544
rect 162400 71324 162452 71330
rect 162400 71266 162452 71272
rect 161860 70366 162072 70394
rect 162136 70366 162348 70394
rect 161676 69902 161704 70366
rect 161664 69896 161716 69902
rect 161664 69838 161716 69844
rect 161572 45008 161624 45014
rect 161572 44950 161624 44956
rect 162044 28422 162072 70366
rect 162032 28416 162084 28422
rect 162032 28358 162084 28364
rect 162320 27130 162348 70366
rect 162308 27124 162360 27130
rect 162308 27066 162360 27072
rect 162412 25770 162440 71266
rect 162492 70236 162544 70242
rect 162492 70178 162544 70184
rect 162504 69902 162532 70178
rect 162492 69896 162544 69902
rect 162492 69838 162544 69844
rect 162400 25764 162452 25770
rect 162400 25706 162452 25712
rect 162504 10470 162532 69838
rect 162492 10464 162544 10470
rect 162492 10406 162544 10412
rect 161388 9172 161440 9178
rect 161388 9114 161440 9120
rect 161296 6384 161348 6390
rect 161296 6326 161348 6332
rect 162596 4962 162624 71538
rect 162688 11898 162716 74990
rect 162676 11892 162728 11898
rect 162676 11834 162728 11840
rect 162780 10402 162808 79591
rect 162872 76702 162900 79727
rect 162952 79698 163004 79704
rect 162964 77926 162992 79698
rect 163228 79688 163280 79694
rect 163226 79656 163228 79665
rect 163280 79656 163282 79665
rect 163562 79642 163590 80036
rect 163654 79676 163682 80036
rect 163746 79966 163774 80036
rect 163734 79960 163786 79966
rect 163734 79902 163786 79908
rect 163838 79898 163866 80036
rect 163930 79937 163958 80036
rect 164022 79966 164050 80036
rect 164114 79966 164142 80036
rect 164010 79960 164062 79966
rect 163916 79928 163972 79937
rect 163826 79892 163878 79898
rect 164010 79902 164062 79908
rect 164102 79960 164154 79966
rect 164102 79902 164154 79908
rect 164206 79898 164234 80036
rect 164298 79898 164326 80036
rect 164390 79937 164418 80036
rect 164482 79966 164510 80036
rect 164470 79960 164522 79966
rect 164376 79928 164432 79937
rect 163916 79863 163972 79872
rect 164194 79892 164246 79898
rect 163826 79834 163878 79840
rect 164194 79834 164246 79840
rect 164286 79892 164338 79898
rect 164470 79902 164522 79908
rect 164376 79863 164432 79872
rect 164286 79834 164338 79840
rect 164102 79824 164154 79830
rect 164422 79792 164478 79801
rect 164154 79772 164188 79778
rect 164102 79766 164188 79772
rect 164114 79750 164188 79766
rect 163654 79648 163728 79676
rect 163044 79620 163096 79626
rect 163226 79591 163282 79600
rect 163320 79620 163372 79626
rect 163044 79562 163096 79568
rect 162952 77920 163004 77926
rect 162952 77862 163004 77868
rect 163056 76786 163084 79562
rect 163136 79552 163188 79558
rect 163136 79494 163188 79500
rect 162964 76758 163084 76786
rect 162860 76696 162912 76702
rect 162860 76638 162912 76644
rect 162860 76492 162912 76498
rect 162860 76434 162912 76440
rect 162872 43450 162900 76434
rect 162964 62082 162992 76758
rect 163044 76696 163096 76702
rect 163044 76638 163096 76644
rect 163056 69834 163084 76638
rect 163148 75750 163176 79494
rect 163240 78402 163268 79591
rect 163320 79562 163372 79568
rect 163516 79614 163590 79642
rect 163228 78396 163280 78402
rect 163228 78338 163280 78344
rect 163332 76129 163360 79562
rect 163516 79257 163544 79614
rect 163596 79484 163648 79490
rect 163596 79426 163648 79432
rect 163502 79248 163558 79257
rect 163502 79183 163558 79192
rect 163412 78464 163464 78470
rect 163412 78406 163464 78412
rect 163318 76120 163374 76129
rect 163318 76055 163374 76064
rect 163136 75744 163188 75750
rect 163136 75686 163188 75692
rect 163424 72962 163452 78406
rect 163516 77858 163544 79183
rect 163504 77852 163556 77858
rect 163504 77794 163556 77800
rect 163504 77444 163556 77450
rect 163504 77386 163556 77392
rect 163412 72956 163464 72962
rect 163412 72898 163464 72904
rect 163516 70394 163544 77386
rect 163608 75886 163636 79426
rect 163700 75993 163728 79648
rect 163778 79656 163834 79665
rect 164160 79642 164188 79750
rect 164332 79756 164384 79762
rect 164574 79744 164602 80036
rect 164666 79812 164694 80036
rect 164758 79937 164786 80036
rect 164850 79966 164878 80036
rect 164942 79966 164970 80036
rect 164838 79960 164890 79966
rect 164744 79928 164800 79937
rect 164838 79902 164890 79908
rect 164930 79960 164982 79966
rect 164930 79902 164982 79908
rect 164744 79863 164800 79872
rect 164666 79801 164740 79812
rect 164666 79792 164754 79801
rect 164666 79784 164698 79792
rect 164422 79727 164478 79736
rect 164332 79698 164384 79704
rect 163778 79591 163780 79600
rect 163832 79591 163834 79600
rect 163872 79620 163924 79626
rect 163780 79562 163832 79568
rect 163872 79562 163924 79568
rect 164068 79614 164188 79642
rect 164238 79656 164294 79665
rect 163686 75984 163742 75993
rect 163686 75919 163742 75928
rect 163596 75880 163648 75886
rect 163596 75822 163648 75828
rect 163688 72956 163740 72962
rect 163688 72898 163740 72904
rect 163516 70366 163636 70394
rect 163044 69828 163096 69834
rect 163044 69770 163096 69776
rect 163608 68814 163636 70366
rect 163596 68808 163648 68814
rect 163596 68750 163648 68756
rect 162952 62076 163004 62082
rect 162952 62018 163004 62024
rect 162860 43444 162912 43450
rect 162860 43386 162912 43392
rect 163700 31278 163728 72898
rect 163792 43518 163820 79562
rect 163884 76922 163912 79562
rect 164068 79529 164096 79614
rect 164238 79591 164240 79600
rect 164292 79591 164294 79600
rect 164240 79562 164292 79568
rect 164054 79520 164110 79529
rect 164054 79455 164110 79464
rect 163964 79280 164016 79286
rect 163964 79222 164016 79228
rect 163976 78946 164004 79222
rect 163964 78940 164016 78946
rect 163964 78882 164016 78888
rect 164068 77518 164096 79455
rect 164148 78396 164200 78402
rect 164148 78338 164200 78344
rect 164056 77512 164108 77518
rect 164056 77454 164108 77460
rect 163884 76894 164096 76922
rect 163872 75880 163924 75886
rect 163872 75822 163924 75828
rect 163884 70394 163912 75822
rect 164068 71505 164096 76894
rect 164054 71496 164110 71505
rect 164054 71431 164110 71440
rect 163884 70366 164004 70394
rect 163872 70032 163924 70038
rect 163872 69974 163924 69980
rect 163884 69834 163912 69974
rect 163872 69828 163924 69834
rect 163872 69770 163924 69776
rect 163780 43512 163832 43518
rect 163780 43454 163832 43460
rect 163884 33998 163912 69770
rect 163872 33992 163924 33998
rect 163872 33934 163924 33940
rect 163688 31272 163740 31278
rect 163688 31214 163740 31220
rect 163976 24274 164004 70366
rect 163964 24268 164016 24274
rect 163964 24210 164016 24216
rect 164068 14550 164096 71431
rect 164160 15978 164188 78338
rect 164252 76498 164280 79562
rect 164240 76492 164292 76498
rect 164240 76434 164292 76440
rect 164240 76220 164292 76226
rect 164240 76162 164292 76168
rect 164252 42294 164280 76162
rect 164344 69970 164372 79698
rect 164436 79558 164464 79727
rect 164528 79716 164602 79744
rect 164698 79727 164754 79736
rect 164928 79792 164984 79801
rect 164928 79727 164930 79736
rect 164424 79552 164476 79558
rect 164424 79494 164476 79500
rect 164424 79348 164476 79354
rect 164424 79290 164476 79296
rect 164436 78606 164464 79290
rect 164424 78600 164476 78606
rect 164424 78542 164476 78548
rect 164528 77330 164556 79716
rect 164712 79676 164740 79727
rect 164982 79727 164984 79736
rect 165034 79744 165062 80036
rect 165126 79812 165154 80036
rect 165218 79966 165246 80036
rect 165206 79960 165258 79966
rect 165310 79937 165338 80036
rect 165206 79902 165258 79908
rect 165296 79928 165352 79937
rect 165296 79863 165352 79872
rect 165252 79824 165304 79830
rect 165126 79784 165200 79812
rect 165034 79716 165108 79744
rect 164930 79698 164982 79704
rect 164620 79648 164740 79676
rect 164792 79688 164844 79694
rect 164620 77586 164648 79648
rect 164792 79630 164844 79636
rect 164700 79552 164752 79558
rect 164804 79529 164832 79630
rect 165080 79626 165108 79716
rect 164884 79620 164936 79626
rect 164884 79562 164936 79568
rect 165068 79620 165120 79626
rect 165068 79562 165120 79568
rect 164700 79494 164752 79500
rect 164790 79520 164846 79529
rect 164608 77580 164660 77586
rect 164608 77522 164660 77528
rect 164712 77450 164740 79494
rect 164790 79455 164846 79464
rect 164700 77444 164752 77450
rect 164700 77386 164752 77392
rect 164528 77302 164740 77330
rect 164608 76084 164660 76090
rect 164608 76026 164660 76032
rect 164516 75948 164568 75954
rect 164516 75890 164568 75896
rect 164424 75812 164476 75818
rect 164424 75754 164476 75760
rect 164332 69964 164384 69970
rect 164332 69906 164384 69912
rect 164436 69766 164464 75754
rect 164528 69902 164556 75890
rect 164516 69896 164568 69902
rect 164516 69838 164568 69844
rect 164620 69834 164648 76026
rect 164712 72962 164740 77302
rect 164896 76090 164924 79562
rect 164976 79552 165028 79558
rect 164976 79494 165028 79500
rect 164988 76129 165016 79494
rect 165068 79484 165120 79490
rect 165068 79426 165120 79432
rect 165080 77625 165108 79426
rect 165066 77616 165122 77625
rect 165066 77551 165122 77560
rect 165068 77444 165120 77450
rect 165068 77386 165120 77392
rect 164974 76120 165030 76129
rect 164884 76084 164936 76090
rect 164974 76055 165030 76064
rect 164884 76026 164936 76032
rect 164792 75132 164844 75138
rect 164792 75074 164844 75080
rect 164700 72956 164752 72962
rect 164700 72898 164752 72904
rect 164608 69828 164660 69834
rect 164608 69770 164660 69776
rect 164424 69760 164476 69766
rect 164424 69702 164476 69708
rect 164804 66978 164832 75074
rect 164976 70168 165028 70174
rect 164976 70110 165028 70116
rect 164988 69970 165016 70110
rect 164976 69964 165028 69970
rect 164976 69906 165028 69912
rect 164792 66972 164844 66978
rect 164792 66914 164844 66920
rect 164240 42288 164292 42294
rect 164240 42230 164292 42236
rect 164988 31210 165016 69906
rect 165080 33930 165108 77386
rect 165172 75954 165200 79784
rect 165252 79766 165304 79772
rect 165264 79257 165292 79766
rect 165402 79744 165430 80036
rect 165494 79898 165522 80036
rect 165482 79892 165534 79898
rect 165482 79834 165534 79840
rect 165586 79778 165614 80036
rect 165678 79971 165706 80036
rect 165664 79962 165720 79971
rect 165664 79897 165720 79906
rect 165770 79830 165798 80036
rect 165758 79824 165810 79830
rect 165586 79750 165660 79778
rect 165862 79812 165890 80036
rect 165954 79966 165982 80036
rect 165942 79960 165994 79966
rect 166046 79937 166074 80036
rect 166138 79966 166166 80036
rect 166230 79966 166258 80036
rect 166322 79966 166350 80036
rect 166414 79966 166442 80036
rect 166506 79966 166534 80036
rect 166126 79960 166178 79966
rect 165942 79902 165994 79908
rect 166032 79928 166088 79937
rect 166126 79902 166178 79908
rect 166218 79960 166270 79966
rect 166218 79902 166270 79908
rect 166310 79960 166362 79966
rect 166310 79902 166362 79908
rect 166402 79960 166454 79966
rect 166402 79902 166454 79908
rect 166494 79960 166546 79966
rect 166598 79937 166626 80036
rect 166494 79902 166546 79908
rect 166584 79928 166640 79937
rect 166032 79863 166088 79872
rect 166584 79863 166640 79872
rect 166080 79824 166132 79830
rect 165862 79801 165936 79812
rect 165862 79792 165950 79801
rect 165862 79784 165894 79792
rect 165758 79766 165810 79772
rect 165402 79716 165476 79744
rect 165344 79620 165396 79626
rect 165344 79562 165396 79568
rect 165250 79248 165306 79257
rect 165250 79183 165306 79192
rect 165264 77790 165292 79183
rect 165252 77784 165304 77790
rect 165252 77726 165304 77732
rect 165160 75948 165212 75954
rect 165160 75890 165212 75896
rect 165356 70394 165384 79562
rect 165448 75818 165476 79716
rect 165632 79676 165660 79750
rect 166598 79812 166626 79863
rect 166080 79766 166132 79772
rect 166552 79784 166626 79812
rect 165894 79727 165950 79736
rect 165804 79688 165856 79694
rect 165526 79656 165582 79665
rect 165632 79648 165752 79676
rect 165526 79591 165582 79600
rect 165436 75812 165488 75818
rect 165436 75754 165488 75760
rect 165436 72956 165488 72962
rect 165436 72898 165488 72904
rect 165264 70366 165384 70394
rect 165160 70032 165212 70038
rect 165160 69974 165212 69980
rect 165172 69834 165200 69974
rect 165160 69828 165212 69834
rect 165160 69770 165212 69776
rect 165068 33924 165120 33930
rect 165068 33866 165120 33872
rect 164976 31204 165028 31210
rect 164976 31146 165028 31152
rect 165172 22914 165200 69770
rect 165264 25702 165292 70366
rect 165344 70100 165396 70106
rect 165344 70042 165396 70048
rect 165356 69902 165384 70042
rect 165344 69896 165396 69902
rect 165344 69838 165396 69844
rect 165252 25696 165304 25702
rect 165252 25638 165304 25644
rect 165160 22908 165212 22914
rect 165160 22850 165212 22856
rect 164884 17264 164936 17270
rect 164884 17206 164936 17212
rect 164148 15972 164200 15978
rect 164148 15914 164200 15920
rect 164056 14544 164108 14550
rect 164056 14486 164108 14492
rect 162768 10396 162820 10402
rect 162768 10338 162820 10344
rect 162584 4956 162636 4962
rect 162584 4898 162636 4904
rect 161294 4856 161350 4865
rect 161294 4791 161350 4800
rect 161308 480 161336 4791
rect 162492 3868 162544 3874
rect 162492 3810 162544 3816
rect 162504 480 162532 3810
rect 163688 3800 163740 3806
rect 163688 3742 163740 3748
rect 163700 480 163728 3742
rect 164516 3732 164568 3738
rect 164516 3674 164568 3680
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164528 354 164556 3674
rect 164896 3602 164924 17206
rect 165356 15910 165384 69838
rect 165344 15904 165396 15910
rect 165344 15846 165396 15852
rect 165448 13190 165476 72898
rect 165540 17474 165568 79591
rect 165620 79484 165672 79490
rect 165620 79426 165672 79432
rect 165528 17468 165580 17474
rect 165528 17410 165580 17416
rect 165436 13184 165488 13190
rect 165436 13126 165488 13132
rect 165632 11830 165660 79426
rect 165724 79286 165752 79648
rect 165804 79630 165856 79636
rect 165712 79280 165764 79286
rect 165712 79222 165764 79228
rect 165710 79112 165766 79121
rect 165710 79047 165766 79056
rect 165724 40866 165752 79047
rect 165816 78674 165844 79630
rect 165988 79552 166040 79558
rect 165988 79494 166040 79500
rect 165896 79280 165948 79286
rect 165896 79222 165948 79228
rect 165804 78668 165856 78674
rect 165804 78610 165856 78616
rect 165908 78520 165936 79222
rect 165816 78492 165936 78520
rect 165816 76226 165844 78492
rect 165896 78396 165948 78402
rect 165896 78338 165948 78344
rect 165804 76220 165856 76226
rect 165804 76162 165856 76168
rect 165804 75812 165856 75818
rect 165804 75754 165856 75760
rect 165816 67590 165844 75754
rect 165908 69902 165936 78338
rect 166000 73098 166028 79494
rect 166092 75818 166120 79766
rect 166172 79756 166224 79762
rect 166172 79698 166224 79704
rect 166448 79756 166500 79762
rect 166448 79698 166500 79704
rect 166184 78402 166212 79698
rect 166356 79620 166408 79626
rect 166356 79562 166408 79568
rect 166172 78396 166224 78402
rect 166172 78338 166224 78344
rect 166172 78260 166224 78266
rect 166172 78202 166224 78208
rect 166080 75812 166132 75818
rect 166080 75754 166132 75760
rect 165988 73092 166040 73098
rect 165988 73034 166040 73040
rect 166184 72554 166212 78202
rect 166264 75744 166316 75750
rect 166264 75686 166316 75692
rect 166172 72548 166224 72554
rect 166172 72490 166224 72496
rect 166276 70394 166304 75686
rect 166368 75410 166396 79562
rect 166460 75993 166488 79698
rect 166446 75984 166502 75993
rect 166446 75919 166502 75928
rect 166356 75404 166408 75410
rect 166356 75346 166408 75352
rect 166276 70366 166396 70394
rect 165896 69896 165948 69902
rect 165896 69838 165948 69844
rect 165804 67584 165856 67590
rect 165804 67526 165856 67532
rect 166368 62014 166396 70366
rect 166356 62008 166408 62014
rect 166356 61950 166408 61956
rect 166552 42226 166580 79784
rect 166690 79778 166718 80036
rect 166782 79898 166810 80036
rect 166874 79898 166902 80036
rect 166966 79937 166994 80036
rect 166952 79928 167008 79937
rect 166770 79892 166822 79898
rect 166770 79834 166822 79840
rect 166862 79892 166914 79898
rect 166952 79863 167008 79872
rect 166862 79834 166914 79840
rect 166690 79750 166764 79778
rect 166632 79688 166684 79694
rect 166630 79656 166632 79665
rect 166736 79676 166764 79750
rect 167058 79744 167086 80036
rect 167150 79937 167178 80036
rect 167242 79966 167270 80036
rect 167230 79960 167282 79966
rect 167136 79928 167192 79937
rect 167230 79902 167282 79908
rect 167334 79903 167362 80036
rect 167136 79863 167192 79872
rect 167320 79894 167376 79903
rect 167320 79829 167376 79838
rect 167426 79778 167454 80036
rect 167518 79937 167546 80036
rect 167504 79928 167560 79937
rect 167504 79863 167560 79872
rect 167426 79750 167500 79778
rect 166920 79716 167086 79744
rect 166684 79656 166686 79665
rect 166736 79648 166856 79676
rect 166630 79591 166686 79600
rect 166644 78577 166672 79591
rect 166724 79552 166776 79558
rect 166724 79494 166776 79500
rect 166630 78568 166686 78577
rect 166630 78503 166686 78512
rect 166736 78146 166764 79494
rect 166644 78118 166764 78146
rect 166644 71194 166672 78118
rect 166722 78024 166778 78033
rect 166722 77959 166778 77968
rect 166632 71188 166684 71194
rect 166632 71130 166684 71136
rect 166632 69896 166684 69902
rect 166632 69838 166684 69844
rect 166540 42220 166592 42226
rect 166540 42162 166592 42168
rect 165712 40860 165764 40866
rect 165712 40802 165764 40808
rect 166644 29782 166672 69838
rect 166736 32502 166764 77959
rect 166828 75993 166856 79648
rect 166814 75984 166870 75993
rect 166814 75919 166870 75928
rect 166920 75818 166948 79716
rect 167090 79656 167146 79665
rect 167000 79620 167052 79626
rect 167274 79656 167330 79665
rect 167090 79591 167146 79600
rect 167184 79620 167236 79626
rect 167000 79562 167052 79568
rect 167012 79257 167040 79562
rect 166998 79248 167054 79257
rect 166998 79183 167054 79192
rect 167012 78402 167040 79183
rect 167000 78396 167052 78402
rect 167000 78338 167052 78344
rect 167104 76106 167132 79591
rect 167274 79591 167330 79600
rect 167184 79562 167236 79568
rect 167196 76702 167224 79562
rect 167184 76696 167236 76702
rect 167184 76638 167236 76644
rect 167012 76078 167132 76106
rect 166908 75812 166960 75818
rect 166908 75754 166960 75760
rect 166908 75404 166960 75410
rect 166908 75346 166960 75352
rect 166920 74526 166948 75346
rect 166908 74520 166960 74526
rect 166908 74462 166960 74468
rect 166816 71188 166868 71194
rect 166816 71130 166868 71136
rect 166724 32496 166776 32502
rect 166724 32438 166776 32444
rect 166632 29776 166684 29782
rect 166632 29718 166684 29724
rect 166828 17406 166856 71130
rect 166816 17400 166868 17406
rect 166816 17342 166868 17348
rect 165620 11824 165672 11830
rect 165620 11766 165672 11772
rect 166920 9110 166948 74462
rect 167012 72894 167040 76078
rect 167092 75948 167144 75954
rect 167092 75890 167144 75896
rect 167000 72888 167052 72894
rect 167000 72830 167052 72836
rect 167000 72344 167052 72350
rect 167000 72286 167052 72292
rect 167012 39438 167040 72286
rect 167104 69018 167132 75890
rect 167184 75812 167236 75818
rect 167184 75754 167236 75760
rect 167196 70378 167224 75754
rect 167184 70372 167236 70378
rect 167184 70314 167236 70320
rect 167288 70310 167316 79591
rect 167472 79529 167500 79750
rect 167610 79744 167638 80036
rect 167702 79966 167730 80036
rect 167794 79971 167822 80036
rect 167690 79960 167742 79966
rect 167690 79902 167742 79908
rect 167780 79962 167836 79971
rect 167780 79897 167836 79906
rect 167610 79716 167776 79744
rect 167550 79656 167606 79665
rect 167550 79591 167606 79600
rect 167458 79520 167514 79529
rect 167458 79455 167514 79464
rect 167368 79212 167420 79218
rect 167368 79154 167420 79160
rect 167380 79121 167408 79154
rect 167366 79112 167422 79121
rect 167366 79047 167422 79056
rect 167472 78334 167500 79455
rect 167564 79121 167592 79591
rect 167550 79112 167606 79121
rect 167550 79047 167606 79056
rect 167460 78328 167512 78334
rect 167460 78270 167512 78276
rect 167644 77376 167696 77382
rect 167644 77318 167696 77324
rect 167656 70394 167684 77318
rect 167748 75954 167776 79716
rect 167886 79608 167914 80036
rect 167978 79812 168006 80036
rect 168070 79937 168098 80036
rect 168056 79928 168112 79937
rect 168056 79863 168112 79872
rect 167978 79784 168052 79812
rect 168024 79676 168052 79784
rect 168162 79744 168190 80036
rect 168254 79971 168282 80036
rect 168240 79962 168296 79971
rect 168346 79966 168374 80036
rect 168438 79966 168466 80036
rect 168530 79966 168558 80036
rect 168240 79897 168296 79906
rect 168334 79960 168386 79966
rect 168334 79902 168386 79908
rect 168426 79960 168478 79966
rect 168426 79902 168478 79908
rect 168518 79960 168570 79966
rect 168518 79902 168570 79908
rect 168288 79824 168340 79830
rect 168288 79766 168340 79772
rect 168424 79826 168480 79835
rect 168622 79830 168650 80036
rect 168162 79716 168236 79744
rect 168024 79665 168144 79676
rect 167840 79580 167914 79608
rect 168010 79656 168144 79665
rect 168066 79648 168144 79656
rect 168010 79591 168066 79600
rect 167736 75948 167788 75954
rect 167736 75890 167788 75896
rect 167840 73166 167868 79580
rect 168012 79552 168064 79558
rect 168010 79520 168012 79529
rect 168064 79520 168066 79529
rect 167932 79478 168010 79506
rect 167828 73160 167880 73166
rect 167828 73102 167880 73108
rect 167656 70366 167776 70394
rect 167276 70304 167328 70310
rect 167276 70246 167328 70252
rect 167092 69012 167144 69018
rect 167092 68954 167144 68960
rect 167000 39432 167052 39438
rect 167000 39374 167052 39380
rect 167000 35216 167052 35222
rect 167000 35158 167052 35164
rect 167012 16574 167040 35158
rect 167748 29850 167776 70366
rect 167828 70304 167880 70310
rect 167828 70246 167880 70252
rect 167840 38078 167868 70246
rect 167828 38072 167880 38078
rect 167828 38014 167880 38020
rect 167932 35358 167960 79478
rect 168010 79455 168066 79464
rect 168116 79404 168144 79648
rect 168024 79376 168144 79404
rect 168024 75206 168052 79376
rect 168104 79008 168156 79014
rect 168104 78950 168156 78956
rect 168012 75200 168064 75206
rect 168012 75142 168064 75148
rect 168012 73160 168064 73166
rect 168012 73102 168064 73108
rect 167920 35352 167972 35358
rect 167920 35294 167972 35300
rect 167736 29844 167788 29850
rect 167736 29786 167788 29792
rect 168024 28354 168052 73102
rect 168116 72350 168144 78950
rect 168208 75993 168236 79716
rect 168300 79014 168328 79766
rect 168424 79761 168480 79770
rect 168610 79824 168662 79830
rect 168714 79812 168742 80036
rect 168806 79937 168834 80036
rect 168898 79966 168926 80036
rect 168886 79960 168938 79966
rect 168792 79928 168848 79937
rect 168886 79902 168938 79908
rect 168990 79898 169018 80036
rect 169082 79966 169110 80036
rect 169174 79971 169202 80036
rect 169070 79960 169122 79966
rect 169070 79902 169122 79908
rect 169160 79962 169216 79971
rect 168792 79863 168848 79872
rect 168978 79892 169030 79898
rect 169160 79897 169216 79906
rect 168978 79834 169030 79840
rect 169116 79824 169168 79830
rect 168714 79784 168788 79812
rect 168610 79766 168662 79772
rect 168760 79778 168788 79784
rect 169022 79792 169078 79801
rect 168438 79676 168466 79761
rect 168760 79750 168834 79778
rect 168438 79648 168512 79676
rect 168378 79520 168434 79529
rect 168378 79455 168434 79464
rect 168288 79008 168340 79014
rect 168288 78950 168340 78956
rect 168286 78704 168342 78713
rect 168286 78639 168342 78648
rect 168194 75984 168250 75993
rect 168194 75919 168250 75928
rect 168104 72344 168156 72350
rect 168104 72286 168156 72292
rect 168300 70394 168328 78639
rect 168104 70372 168156 70378
rect 168104 70314 168156 70320
rect 168208 70366 168328 70394
rect 168012 28348 168064 28354
rect 168012 28290 168064 28296
rect 168116 17338 168144 70314
rect 168208 22846 168236 70366
rect 168288 69012 168340 69018
rect 168288 68954 168340 68960
rect 168196 22840 168248 22846
rect 168196 22782 168248 22788
rect 168104 17332 168156 17338
rect 168104 17274 168156 17280
rect 167012 16546 167224 16574
rect 166908 9104 166960 9110
rect 166908 9046 166960 9052
rect 166080 3732 166132 3738
rect 166080 3674 166132 3680
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 166092 480 166120 3674
rect 167196 480 167224 16546
rect 168300 7682 168328 68954
rect 168392 46306 168420 79455
rect 168380 46300 168432 46306
rect 168380 46242 168432 46248
rect 168484 39506 168512 79648
rect 168806 79642 168834 79750
rect 169116 79766 169168 79772
rect 169022 79727 169078 79736
rect 169036 79642 169064 79727
rect 168564 79620 168616 79626
rect 168564 79562 168616 79568
rect 168656 79620 168708 79626
rect 168656 79562 168708 79568
rect 168760 79614 168834 79642
rect 168944 79614 169064 79642
rect 168576 77761 168604 79562
rect 168562 77752 168618 77761
rect 168562 77687 168618 77696
rect 168564 76492 168616 76498
rect 168564 76434 168616 76440
rect 168576 53786 168604 76434
rect 168668 55214 168696 79562
rect 168760 76498 168788 79614
rect 168840 79552 168892 79558
rect 168840 79494 168892 79500
rect 168748 76492 168800 76498
rect 168748 76434 168800 76440
rect 168852 76430 168880 79494
rect 168944 78826 168972 79614
rect 169022 79248 169078 79257
rect 169022 79183 169078 79192
rect 169036 78946 169064 79183
rect 169024 78940 169076 78946
rect 169024 78882 169076 78888
rect 168944 78798 169064 78826
rect 168930 78296 168986 78305
rect 168930 78231 168986 78240
rect 168840 76424 168892 76430
rect 168840 76366 168892 76372
rect 168944 75914 168972 78231
rect 169036 76498 169064 78798
rect 169128 76945 169156 79766
rect 169266 79744 169294 80036
rect 169358 79898 169386 80036
rect 169450 79971 169478 80036
rect 169436 79962 169492 79971
rect 169346 79892 169398 79898
rect 169436 79897 169492 79906
rect 169346 79834 169398 79840
rect 169542 79812 169570 80036
rect 169634 79898 169662 80036
rect 169726 79966 169754 80036
rect 169818 79966 169846 80036
rect 169714 79960 169766 79966
rect 169714 79902 169766 79908
rect 169806 79960 169858 79966
rect 169806 79902 169858 79908
rect 169910 79898 169938 80036
rect 170002 79966 170030 80036
rect 170094 79971 170122 80036
rect 169990 79960 170042 79966
rect 169990 79902 170042 79908
rect 170080 79962 170136 79971
rect 169622 79892 169674 79898
rect 169622 79834 169674 79840
rect 169898 79892 169950 79898
rect 170080 79897 170136 79906
rect 169898 79834 169950 79840
rect 169496 79784 169570 79812
rect 169266 79716 169340 79744
rect 169208 79620 169260 79626
rect 169208 79562 169260 79568
rect 169220 79529 169248 79562
rect 169206 79520 169262 79529
rect 169206 79455 169262 79464
rect 169220 78946 169248 79455
rect 169208 78940 169260 78946
rect 169312 78928 169340 79716
rect 169390 79656 169446 79665
rect 169390 79591 169392 79600
rect 169444 79591 169446 79600
rect 169392 79562 169444 79568
rect 169392 79484 169444 79490
rect 169496 79472 169524 79784
rect 169852 79756 169904 79762
rect 170186 79744 170214 80036
rect 170278 79966 170306 80036
rect 170266 79960 170318 79966
rect 170266 79902 170318 79908
rect 170370 79898 170398 80036
rect 170462 79937 170490 80036
rect 170554 79966 170582 80036
rect 170542 79960 170594 79966
rect 170448 79928 170504 79937
rect 170358 79892 170410 79898
rect 170542 79902 170594 79908
rect 170448 79863 170504 79872
rect 170358 79834 170410 79840
rect 170646 79812 170674 80036
rect 170738 79966 170766 80036
rect 170726 79960 170778 79966
rect 170726 79902 170778 79908
rect 170646 79784 170720 79812
rect 170186 79716 170536 79744
rect 169852 79698 169904 79704
rect 169668 79620 169720 79626
rect 169668 79562 169720 79568
rect 169496 79444 169616 79472
rect 169392 79426 169444 79432
rect 169404 79393 169432 79426
rect 169390 79384 169446 79393
rect 169446 79342 169524 79370
rect 169390 79319 169446 79328
rect 169312 78900 169432 78928
rect 169208 78882 169260 78888
rect 169114 76936 169170 76945
rect 169114 76871 169170 76880
rect 169116 76696 169168 76702
rect 169116 76638 169168 76644
rect 169024 76492 169076 76498
rect 169024 76434 169076 76440
rect 168852 75886 168972 75914
rect 168748 75132 168800 75138
rect 168748 75074 168800 75080
rect 168760 57934 168788 75074
rect 168852 64870 168880 75886
rect 169128 69834 169156 76638
rect 169208 76424 169260 76430
rect 169208 76366 169260 76372
rect 169116 69828 169168 69834
rect 169116 69770 169168 69776
rect 168840 64864 168892 64870
rect 168840 64806 168892 64812
rect 168748 57928 168800 57934
rect 168748 57870 168800 57876
rect 168656 55208 168708 55214
rect 168656 55150 168708 55156
rect 168564 53780 168616 53786
rect 168564 53722 168616 53728
rect 169220 52426 169248 76366
rect 169404 75914 169432 78900
rect 169496 77994 169524 79342
rect 169484 77988 169536 77994
rect 169484 77930 169536 77936
rect 169312 75886 169432 75914
rect 169588 75914 169616 79444
rect 169680 78606 169708 79562
rect 169760 79552 169812 79558
rect 169760 79494 169812 79500
rect 169772 79121 169800 79494
rect 169864 79472 169892 79698
rect 170036 79688 170088 79694
rect 170036 79630 170088 79636
rect 169864 79444 169984 79472
rect 169758 79112 169814 79121
rect 169814 79070 169892 79098
rect 169758 79047 169814 79056
rect 169668 78600 169720 78606
rect 169668 78542 169720 78548
rect 169864 78266 169892 79070
rect 169852 78260 169904 78266
rect 169852 78202 169904 78208
rect 169760 77988 169812 77994
rect 169760 77930 169812 77936
rect 169588 75886 169708 75914
rect 169312 75138 169340 75886
rect 169300 75132 169352 75138
rect 169300 75074 169352 75080
rect 169680 71534 169708 75886
rect 169668 71528 169720 71534
rect 169668 71470 169720 71476
rect 169208 52420 169260 52426
rect 169208 52362 169260 52368
rect 169024 51876 169076 51882
rect 169024 51818 169076 51824
rect 168564 47592 168616 47598
rect 168564 47534 168616 47540
rect 168472 39500 168524 39506
rect 168472 39442 168524 39448
rect 168576 16574 168604 47534
rect 168576 16546 168972 16574
rect 168288 7676 168340 7682
rect 168288 7618 168340 7624
rect 168380 3596 168432 3602
rect 168380 3538 168432 3544
rect 168392 480 168420 3538
rect 168944 3482 168972 16546
rect 169036 4146 169064 51818
rect 169680 17270 169708 71470
rect 169668 17264 169720 17270
rect 169668 17206 169720 17212
rect 169772 6322 169800 77930
rect 169852 77716 169904 77722
rect 169852 77658 169904 77664
rect 169864 31074 169892 77658
rect 169956 77382 169984 79444
rect 170048 78470 170076 79630
rect 170220 79620 170272 79626
rect 170220 79562 170272 79568
rect 170036 78464 170088 78470
rect 170036 78406 170088 78412
rect 169944 77376 169996 77382
rect 169944 77318 169996 77324
rect 170232 76906 170260 79562
rect 170312 79552 170364 79558
rect 170312 79494 170364 79500
rect 170404 79552 170456 79558
rect 170404 79494 170456 79500
rect 170324 79393 170352 79494
rect 170310 79384 170366 79393
rect 170310 79319 170366 79328
rect 170312 78804 170364 78810
rect 170312 78746 170364 78752
rect 170324 78538 170352 78746
rect 170312 78532 170364 78538
rect 170312 78474 170364 78480
rect 170220 76900 170272 76906
rect 170220 76842 170272 76848
rect 170218 76528 170274 76537
rect 170218 76463 170274 76472
rect 170232 70394 170260 76463
rect 170416 75750 170444 79494
rect 170508 79121 170536 79716
rect 170494 79112 170550 79121
rect 170494 79047 170550 79056
rect 170494 78976 170550 78985
rect 170494 78911 170550 78920
rect 170404 75744 170456 75750
rect 170404 75686 170456 75692
rect 170232 70366 170444 70394
rect 169852 31068 169904 31074
rect 169852 31010 169904 31016
rect 169760 6316 169812 6322
rect 169760 6258 169812 6264
rect 170416 4894 170444 70366
rect 170508 58682 170536 78911
rect 170692 77466 170720 79784
rect 170830 79778 170858 80036
rect 170922 79898 170950 80036
rect 170910 79892 170962 79898
rect 170910 79834 170962 79840
rect 171014 79801 171042 80036
rect 171106 79966 171134 80036
rect 171198 79966 171226 80036
rect 171094 79960 171146 79966
rect 171094 79902 171146 79908
rect 171186 79960 171238 79966
rect 171290 79937 171318 80036
rect 171382 79966 171410 80036
rect 171370 79960 171422 79966
rect 171186 79902 171238 79908
rect 171276 79928 171332 79937
rect 171370 79902 171422 79908
rect 171276 79863 171332 79872
rect 171324 79824 171376 79830
rect 170784 79750 170858 79778
rect 171000 79792 171056 79801
rect 170784 77625 170812 79750
rect 171474 79812 171502 80036
rect 171566 79937 171594 80036
rect 171552 79928 171608 79937
rect 171552 79863 171608 79872
rect 171658 79812 171686 80036
rect 171750 79966 171778 80036
rect 171738 79960 171790 79966
rect 171738 79902 171790 79908
rect 171474 79784 171548 79812
rect 171324 79766 171376 79772
rect 171000 79727 171056 79736
rect 171232 79756 171284 79762
rect 171232 79698 171284 79704
rect 170864 79688 170916 79694
rect 170862 79656 170864 79665
rect 171048 79688 171100 79694
rect 170916 79656 170918 79665
rect 170918 79614 170996 79642
rect 171048 79630 171100 79636
rect 170862 79591 170918 79600
rect 170864 78940 170916 78946
rect 170864 78882 170916 78888
rect 170876 78266 170904 78882
rect 170864 78260 170916 78266
rect 170864 78202 170916 78208
rect 170770 77616 170826 77625
rect 170770 77551 170826 77560
rect 170692 77438 170904 77466
rect 170680 77376 170732 77382
rect 170680 77318 170732 77324
rect 170588 76900 170640 76906
rect 170588 76842 170640 76848
rect 170496 58676 170548 58682
rect 170496 58618 170548 58624
rect 170600 47666 170628 76842
rect 170692 76838 170720 77318
rect 170680 76832 170732 76838
rect 170680 76774 170732 76780
rect 170588 47660 170640 47666
rect 170588 47602 170640 47608
rect 170692 38010 170720 76774
rect 170876 76702 170904 77438
rect 170864 76696 170916 76702
rect 170770 76664 170826 76673
rect 170864 76638 170916 76644
rect 170770 76599 170826 76608
rect 170680 38004 170732 38010
rect 170680 37946 170732 37952
rect 170784 36650 170812 76599
rect 170772 36644 170824 36650
rect 170772 36586 170824 36592
rect 170876 33862 170904 76638
rect 170864 33856 170916 33862
rect 170864 33798 170916 33804
rect 170968 10334 170996 79614
rect 171060 79529 171088 79630
rect 171140 79620 171192 79626
rect 171140 79562 171192 79568
rect 171046 79520 171102 79529
rect 171046 79455 171102 79464
rect 171152 77722 171180 79562
rect 171244 78985 171272 79698
rect 171230 78976 171286 78985
rect 171230 78911 171286 78920
rect 171140 77716 171192 77722
rect 171140 77658 171192 77664
rect 171048 75744 171100 75750
rect 171048 75686 171100 75692
rect 171060 54534 171088 75686
rect 171244 70394 171272 78911
rect 171336 78033 171364 79766
rect 171416 79688 171468 79694
rect 171416 79630 171468 79636
rect 171322 78024 171378 78033
rect 171322 77959 171378 77968
rect 171428 75818 171456 79630
rect 171520 79257 171548 79784
rect 171612 79784 171686 79812
rect 171506 79248 171562 79257
rect 171506 79183 171562 79192
rect 171508 78940 171560 78946
rect 171508 78882 171560 78888
rect 171416 75812 171468 75818
rect 171416 75754 171468 75760
rect 171520 74390 171548 78882
rect 171612 76537 171640 79784
rect 171842 79744 171870 80036
rect 171934 79812 171962 80036
rect 172026 79966 172054 80036
rect 172014 79960 172066 79966
rect 172118 79937 172146 80036
rect 172014 79902 172066 79908
rect 172104 79928 172160 79937
rect 172104 79863 172160 79872
rect 172060 79824 172112 79830
rect 171934 79784 172008 79812
rect 171842 79716 171916 79744
rect 171888 79665 171916 79716
rect 171874 79656 171930 79665
rect 171874 79591 171930 79600
rect 171690 79520 171746 79529
rect 171690 79455 171746 79464
rect 171704 79422 171732 79455
rect 171692 79416 171744 79422
rect 171692 79358 171744 79364
rect 171690 79248 171746 79257
rect 171690 79183 171746 79192
rect 171704 77294 171732 79183
rect 171888 78538 171916 79591
rect 171876 78532 171928 78538
rect 171876 78474 171928 78480
rect 171874 78296 171930 78305
rect 171874 78231 171930 78240
rect 171704 77266 171824 77294
rect 171598 76528 171654 76537
rect 171598 76463 171654 76472
rect 171508 74384 171560 74390
rect 171508 74326 171560 74332
rect 171244 70366 171364 70394
rect 171048 54528 171100 54534
rect 171048 54470 171100 54476
rect 171336 42158 171364 70366
rect 171324 42152 171376 42158
rect 171324 42094 171376 42100
rect 171796 35290 171824 77266
rect 171784 35284 171836 35290
rect 171784 35226 171836 35232
rect 171782 27024 171838 27033
rect 171782 26959 171838 26968
rect 170956 10328 171008 10334
rect 170956 10270 171008 10276
rect 170404 4888 170456 4894
rect 170404 4830 170456 4836
rect 169024 4140 169076 4146
rect 169024 4082 169076 4088
rect 170772 3936 170824 3942
rect 170772 3878 170824 3884
rect 168944 3454 169616 3482
rect 169588 480 169616 3454
rect 170784 480 170812 3878
rect 171796 3194 171824 26959
rect 171888 14482 171916 78231
rect 171980 77897 172008 79784
rect 172210 79812 172238 80036
rect 172302 79937 172330 80036
rect 172394 79966 172422 80036
rect 172382 79960 172434 79966
rect 172288 79928 172344 79937
rect 172382 79902 172434 79908
rect 172288 79863 172344 79872
rect 172336 79824 172388 79830
rect 172210 79784 172284 79812
rect 172060 79766 172112 79772
rect 172072 79608 172100 79766
rect 172072 79580 172192 79608
rect 172058 79520 172114 79529
rect 172058 79455 172114 79464
rect 171966 77888 172022 77897
rect 171966 77823 172022 77832
rect 172072 77772 172100 79455
rect 172164 78946 172192 79580
rect 172256 78985 172284 79784
rect 172336 79766 172388 79772
rect 172348 79257 172376 79766
rect 172486 79744 172514 80036
rect 172440 79716 172514 79744
rect 172578 79744 172606 80036
rect 172670 79812 172698 80036
rect 172762 79971 172790 80036
rect 172748 79962 172804 79971
rect 172854 79966 172882 80036
rect 172946 79971 172974 80036
rect 172748 79897 172804 79906
rect 172842 79960 172894 79966
rect 172842 79902 172894 79908
rect 172932 79962 172988 79971
rect 173038 79966 173066 80036
rect 172932 79897 172988 79906
rect 173026 79960 173078 79966
rect 173026 79902 173078 79908
rect 172980 79824 173032 79830
rect 172670 79784 172744 79812
rect 172578 79716 172652 79744
rect 172334 79248 172390 79257
rect 172334 79183 172390 79192
rect 172242 78976 172298 78985
rect 172152 78940 172204 78946
rect 172242 78911 172298 78920
rect 172152 78882 172204 78888
rect 172244 78532 172296 78538
rect 172244 78474 172296 78480
rect 171980 77744 172100 77772
rect 171980 76362 172008 77744
rect 172058 77616 172114 77625
rect 172058 77551 172114 77560
rect 171968 76356 172020 76362
rect 171968 76298 172020 76304
rect 171980 75954 172008 76298
rect 171968 75948 172020 75954
rect 171968 75890 172020 75896
rect 171968 75812 172020 75818
rect 171968 75754 172020 75760
rect 171980 28286 172008 75754
rect 171968 28280 172020 28286
rect 171968 28222 172020 28228
rect 171876 14476 171928 14482
rect 171876 14418 171928 14424
rect 172072 13122 172100 77551
rect 172152 75948 172204 75954
rect 172152 75890 172204 75896
rect 172164 75154 172192 75890
rect 172256 75342 172284 78474
rect 172244 75336 172296 75342
rect 172244 75278 172296 75284
rect 172348 75274 172376 79183
rect 172440 78577 172468 79716
rect 172624 79608 172652 79716
rect 172532 79580 172652 79608
rect 172426 78568 172482 78577
rect 172426 78503 172482 78512
rect 172336 75268 172388 75274
rect 172336 75210 172388 75216
rect 172164 75126 172284 75154
rect 172152 74384 172204 74390
rect 172152 74326 172204 74332
rect 172164 73710 172192 74326
rect 172152 73704 172204 73710
rect 172152 73646 172204 73652
rect 172164 26994 172192 73646
rect 172152 26988 172204 26994
rect 172152 26930 172204 26936
rect 172256 25634 172284 75126
rect 172532 74322 172560 79580
rect 172716 79506 172744 79784
rect 173130 79778 173158 80036
rect 173222 79966 173250 80036
rect 173314 79966 173342 80036
rect 173406 79966 173434 80036
rect 173210 79960 173262 79966
rect 173210 79902 173262 79908
rect 173302 79960 173354 79966
rect 173302 79902 173354 79908
rect 173394 79960 173446 79966
rect 173498 79937 173526 80036
rect 173394 79902 173446 79908
rect 173484 79928 173540 79937
rect 173590 79898 173618 80036
rect 173682 79966 173710 80036
rect 173774 79966 173802 80036
rect 173866 79971 173894 80036
rect 173670 79960 173722 79966
rect 173670 79902 173722 79908
rect 173762 79960 173814 79966
rect 173762 79902 173814 79908
rect 173852 79962 173908 79971
rect 173958 79966 173986 80036
rect 173484 79863 173540 79872
rect 173578 79892 173630 79898
rect 173852 79897 173908 79906
rect 173946 79960 173998 79966
rect 173946 79902 173998 79908
rect 172980 79766 173032 79772
rect 172796 79756 172848 79762
rect 172796 79698 172848 79704
rect 172808 79608 172836 79698
rect 172808 79580 172928 79608
rect 172716 79478 172790 79506
rect 172762 79472 172790 79478
rect 172762 79444 172836 79472
rect 172612 78940 172664 78946
rect 172612 78882 172664 78888
rect 172624 78810 172652 78882
rect 172612 78804 172664 78810
rect 172612 78746 172664 78752
rect 172808 77246 172836 79444
rect 172796 77240 172848 77246
rect 172796 77182 172848 77188
rect 172704 76084 172756 76090
rect 172704 76026 172756 76032
rect 172520 74316 172572 74322
rect 172520 74258 172572 74264
rect 172520 73772 172572 73778
rect 172520 73714 172572 73720
rect 172532 44946 172560 73714
rect 172716 61878 172744 76026
rect 172900 74390 172928 79580
rect 172992 75410 173020 79766
rect 173084 79750 173158 79778
rect 173256 79824 173308 79830
rect 173256 79766 173308 79772
rect 173348 79824 173400 79830
rect 173348 79766 173400 79772
rect 173084 79257 173112 79750
rect 173268 79665 173296 79766
rect 173254 79656 173310 79665
rect 173254 79591 173310 79600
rect 173254 79520 173310 79529
rect 173254 79455 173310 79464
rect 173070 79248 173126 79257
rect 173070 79183 173126 79192
rect 172980 75404 173032 75410
rect 172980 75346 173032 75352
rect 172888 74384 172940 74390
rect 172888 74326 172940 74332
rect 173084 70394 173112 79183
rect 173164 79076 173216 79082
rect 173164 79018 173216 79024
rect 173176 78810 173204 79018
rect 173164 78804 173216 78810
rect 173164 78746 173216 78752
rect 173084 70366 173204 70394
rect 172704 61872 172756 61878
rect 172704 61814 172756 61820
rect 172520 44940 172572 44946
rect 172520 44882 172572 44888
rect 172244 25628 172296 25634
rect 172244 25570 172296 25576
rect 173176 24206 173204 70366
rect 173268 25566 173296 79455
rect 173360 79121 173388 79766
rect 173498 79744 173526 79863
rect 173578 79834 173630 79840
rect 173716 79824 173768 79830
rect 173716 79766 173768 79772
rect 173624 79756 173676 79762
rect 173498 79716 173572 79744
rect 173346 79112 173402 79121
rect 173346 79047 173402 79056
rect 173360 73778 173388 79047
rect 173544 75970 173572 79716
rect 173624 79698 173676 79704
rect 173636 76090 173664 79698
rect 173728 79529 173756 79766
rect 173808 79756 173860 79762
rect 174050 79744 174078 80036
rect 173808 79698 173860 79704
rect 174004 79716 174078 79744
rect 173714 79520 173770 79529
rect 173714 79455 173770 79464
rect 173820 79200 173848 79698
rect 173900 79688 173952 79694
rect 173900 79630 173952 79636
rect 173728 79172 173848 79200
rect 173728 78656 173756 79172
rect 173808 79076 173860 79082
rect 173808 79018 173860 79024
rect 173820 78810 173848 79018
rect 173808 78804 173860 78810
rect 173808 78746 173860 78752
rect 173728 78628 173848 78656
rect 173714 78568 173770 78577
rect 173714 78503 173770 78512
rect 173624 76084 173676 76090
rect 173624 76026 173676 76032
rect 173544 75942 173664 75970
rect 173532 74384 173584 74390
rect 173532 74326 173584 74332
rect 173440 74316 173492 74322
rect 173440 74258 173492 74264
rect 173348 73772 173400 73778
rect 173348 73714 173400 73720
rect 173452 40798 173480 74258
rect 173440 40792 173492 40798
rect 173440 40734 173492 40740
rect 173544 39370 173572 74326
rect 173636 42090 173664 75942
rect 173624 42084 173676 42090
rect 173624 42026 173676 42032
rect 173532 39364 173584 39370
rect 173532 39306 173584 39312
rect 173728 26926 173756 78503
rect 173820 75993 173848 78628
rect 173806 75984 173862 75993
rect 173806 75919 173862 75928
rect 173912 74361 173940 79630
rect 174004 78928 174032 79716
rect 174142 79676 174170 80036
rect 174234 79898 174262 80036
rect 174326 79937 174354 80036
rect 174418 79966 174446 80036
rect 174406 79960 174458 79966
rect 174312 79928 174368 79937
rect 174222 79892 174274 79898
rect 174406 79902 174458 79908
rect 174510 79898 174538 80036
rect 174602 79966 174630 80036
rect 174694 79966 174722 80036
rect 174786 79966 174814 80036
rect 174590 79960 174642 79966
rect 174590 79902 174642 79908
rect 174682 79960 174734 79966
rect 174682 79902 174734 79908
rect 174774 79960 174826 79966
rect 174774 79902 174826 79908
rect 174312 79863 174368 79872
rect 174498 79892 174550 79898
rect 174222 79834 174274 79840
rect 174498 79834 174550 79840
rect 174878 79830 174906 80036
rect 174970 79898 174998 80036
rect 175062 79898 175090 80036
rect 174958 79892 175010 79898
rect 174958 79834 175010 79840
rect 175050 79892 175102 79898
rect 175050 79834 175102 79840
rect 174360 79824 174412 79830
rect 174728 79824 174780 79830
rect 174360 79766 174412 79772
rect 174542 79792 174598 79801
rect 174096 79648 174170 79676
rect 174096 79529 174124 79648
rect 174082 79520 174138 79529
rect 174082 79455 174138 79464
rect 174176 79484 174228 79490
rect 174176 79426 174228 79432
rect 174004 78900 174124 78928
rect 173992 78804 174044 78810
rect 173992 78746 174044 78752
rect 174004 78062 174032 78746
rect 173992 78056 174044 78062
rect 173992 77998 174044 78004
rect 174096 75721 174124 78900
rect 174188 78062 174216 79426
rect 174372 79354 174400 79766
rect 174598 79762 174676 79778
rect 174728 79766 174780 79772
rect 174866 79824 174918 79830
rect 175154 79801 175182 80036
rect 175246 79937 175274 80036
rect 175232 79928 175288 79937
rect 175232 79863 175288 79872
rect 174866 79766 174918 79772
rect 175140 79792 175196 79801
rect 174598 79756 174688 79762
rect 174598 79750 174636 79756
rect 174542 79727 174598 79736
rect 174636 79698 174688 79704
rect 174544 79688 174596 79694
rect 174544 79630 174596 79636
rect 174360 79348 174412 79354
rect 174360 79290 174412 79296
rect 174176 78056 174228 78062
rect 174176 77998 174228 78004
rect 174082 75712 174138 75721
rect 174082 75647 174138 75656
rect 173898 74352 173954 74361
rect 173898 74287 173954 74296
rect 174372 69014 174400 79290
rect 174556 75449 174584 79630
rect 174542 75440 174598 75449
rect 174542 75375 174598 75384
rect 174004 68986 174400 69014
rect 174004 64874 174032 68986
rect 173912 64846 174032 64874
rect 173716 26920 173768 26926
rect 173716 26862 173768 26868
rect 173256 25560 173308 25566
rect 173256 25502 173308 25508
rect 173164 24200 173216 24206
rect 173164 24142 173216 24148
rect 173256 24132 173308 24138
rect 173256 24074 173308 24080
rect 172060 13116 172112 13122
rect 172060 13058 172112 13064
rect 173164 4140 173216 4146
rect 173164 4082 173216 4088
rect 171968 3664 172020 3670
rect 171968 3606 172020 3612
rect 171784 3188 171836 3194
rect 171784 3130 171836 3136
rect 171980 480 172008 3606
rect 173176 480 173204 4082
rect 173268 3602 173296 24074
rect 173912 4826 173940 64846
rect 174648 44878 174676 79698
rect 174740 75585 174768 79766
rect 175004 79756 175056 79762
rect 175140 79727 175196 79736
rect 175338 79744 175366 80036
rect 175430 79937 175458 80036
rect 175522 79966 175550 80036
rect 175510 79960 175562 79966
rect 175416 79928 175472 79937
rect 175510 79902 175562 79908
rect 175416 79863 175472 79872
rect 175614 79830 175642 80036
rect 175706 79830 175734 80036
rect 175798 79937 175826 80036
rect 175784 79928 175840 79937
rect 175784 79863 175840 79872
rect 175464 79824 175516 79830
rect 175464 79766 175516 79772
rect 175602 79824 175654 79830
rect 175602 79766 175654 79772
rect 175694 79824 175746 79830
rect 175890 79778 175918 80036
rect 175982 79966 176010 80036
rect 175970 79960 176022 79966
rect 175970 79902 176022 79908
rect 175694 79766 175746 79772
rect 175338 79716 175412 79744
rect 175004 79698 175056 79704
rect 174820 79688 174872 79694
rect 174818 79656 174820 79665
rect 174872 79656 174874 79665
rect 174818 79591 174874 79600
rect 174832 78656 174860 79591
rect 174832 78628 174952 78656
rect 174818 78568 174874 78577
rect 174818 78503 174874 78512
rect 174726 75576 174782 75585
rect 174726 75511 174782 75520
rect 174726 75440 174782 75449
rect 174726 75375 174782 75384
rect 174636 44872 174688 44878
rect 174636 44814 174688 44820
rect 174740 37942 174768 75375
rect 174728 37936 174780 37942
rect 174728 37878 174780 37884
rect 174832 32434 174860 78503
rect 174924 76786 174952 78628
rect 175016 76945 175044 79698
rect 175096 79688 175148 79694
rect 175096 79630 175148 79636
rect 175278 79656 175334 79665
rect 175108 77081 175136 79630
rect 175278 79591 175280 79600
rect 175332 79591 175334 79600
rect 175280 79562 175332 79568
rect 175186 79520 175242 79529
rect 175186 79455 175242 79464
rect 175200 78305 175228 79455
rect 175186 78296 175242 78305
rect 175186 78231 175242 78240
rect 175094 77072 175150 77081
rect 175094 77007 175150 77016
rect 175002 76936 175058 76945
rect 175002 76871 175058 76880
rect 174924 76758 175044 76786
rect 174910 74352 174966 74361
rect 174910 74287 174966 74296
rect 174820 32428 174872 32434
rect 174820 32370 174872 32376
rect 174924 22778 174952 74287
rect 175016 24138 175044 76758
rect 175004 24132 175056 24138
rect 175004 24074 175056 24080
rect 174912 22772 174964 22778
rect 174912 22714 174964 22720
rect 175108 11762 175136 77007
rect 175186 73944 175242 73953
rect 175186 73879 175242 73888
rect 175096 11756 175148 11762
rect 175096 11698 175148 11704
rect 175200 7614 175228 73879
rect 175292 49026 175320 79562
rect 175384 79558 175412 79716
rect 175372 79552 175424 79558
rect 175372 79494 175424 79500
rect 175476 73953 175504 79766
rect 175844 79750 175918 79778
rect 175648 79688 175700 79694
rect 175844 79642 175872 79750
rect 176074 79744 176102 80036
rect 176166 79898 176194 80036
rect 176258 79898 176286 80036
rect 176350 79937 176378 80036
rect 176336 79928 176392 79937
rect 176154 79892 176206 79898
rect 176154 79834 176206 79840
rect 176246 79892 176298 79898
rect 176336 79863 176392 79872
rect 176246 79834 176298 79840
rect 176442 79830 176470 80036
rect 176430 79824 176482 79830
rect 176028 79716 176102 79744
rect 176198 79792 176254 79801
rect 176534 79801 176562 80036
rect 176430 79766 176482 79772
rect 176520 79792 176576 79801
rect 176198 79727 176200 79736
rect 175648 79630 175700 79636
rect 175462 73944 175518 73953
rect 175462 73879 175518 73888
rect 175660 72865 175688 79630
rect 175752 79614 175872 79642
rect 175924 79688 175976 79694
rect 175924 79630 175976 79636
rect 175752 78985 175780 79614
rect 175832 79552 175884 79558
rect 175936 79529 175964 79630
rect 175832 79494 175884 79500
rect 175922 79520 175978 79529
rect 175738 78976 175794 78985
rect 175738 78911 175794 78920
rect 175646 72856 175702 72865
rect 175646 72791 175702 72800
rect 175752 69014 175780 78911
rect 175844 74594 175872 79494
rect 175922 79455 175978 79464
rect 175832 74588 175884 74594
rect 175832 74530 175884 74536
rect 175936 72146 175964 79455
rect 176028 78169 176056 79716
rect 176252 79727 176254 79736
rect 176292 79756 176344 79762
rect 176200 79698 176252 79704
rect 176520 79727 176576 79736
rect 176292 79698 176344 79704
rect 176106 79656 176162 79665
rect 176106 79591 176108 79600
rect 176160 79591 176162 79600
rect 176108 79562 176160 79568
rect 176014 78160 176070 78169
rect 176014 78095 176070 78104
rect 176120 78044 176148 79562
rect 176028 78016 176148 78044
rect 175924 72140 175976 72146
rect 175924 72082 175976 72088
rect 176028 70394 176056 78016
rect 176108 74588 176160 74594
rect 176108 74530 176160 74536
rect 176120 72350 176148 74530
rect 176108 72344 176160 72350
rect 176108 72286 176160 72292
rect 175384 68986 175780 69014
rect 175844 70366 176056 70394
rect 175280 49020 175332 49026
rect 175280 48962 175332 48968
rect 175384 29646 175412 68986
rect 175372 29640 175424 29646
rect 175372 29582 175424 29588
rect 175188 7608 175240 7614
rect 175188 7550 175240 7556
rect 175844 6186 175872 70366
rect 176120 36582 176148 72286
rect 176212 40730 176240 79698
rect 176304 77217 176332 79698
rect 176384 79688 176436 79694
rect 176384 79630 176436 79636
rect 176396 77382 176424 79630
rect 176534 79608 176562 79727
rect 176626 79676 176654 80036
rect 176718 79830 176746 80036
rect 176810 79898 176838 80036
rect 176798 79892 176850 79898
rect 176798 79834 176850 79840
rect 176706 79824 176758 79830
rect 176706 79766 176758 79772
rect 176902 79744 176930 80036
rect 176994 79812 177022 80036
rect 177086 79966 177114 80036
rect 177074 79960 177126 79966
rect 177074 79902 177126 79908
rect 176994 79784 177068 79812
rect 176902 79716 176976 79744
rect 176626 79648 176700 79676
rect 176672 79642 176700 79648
rect 176672 79614 176884 79642
rect 176488 79580 176562 79608
rect 176384 77376 176436 77382
rect 176384 77318 176436 77324
rect 176290 77208 176346 77217
rect 176290 77143 176346 77152
rect 176488 75914 176516 79580
rect 176752 79552 176804 79558
rect 176658 79520 176714 79529
rect 176752 79494 176804 79500
rect 176658 79455 176714 79464
rect 176396 75886 176516 75914
rect 176292 72140 176344 72146
rect 176292 72082 176344 72088
rect 176200 40724 176252 40730
rect 176200 40666 176252 40672
rect 176108 36576 176160 36582
rect 176108 36518 176160 36524
rect 176304 18766 176332 72082
rect 176292 18760 176344 18766
rect 176292 18702 176344 18708
rect 176396 18698 176424 75886
rect 176566 75576 176622 75585
rect 176566 75511 176622 75520
rect 176474 72856 176530 72865
rect 176474 72791 176530 72800
rect 176384 18692 176436 18698
rect 176384 18634 176436 18640
rect 176488 9042 176516 72791
rect 176476 9036 176528 9042
rect 176476 8978 176528 8984
rect 176580 6254 176608 75511
rect 176672 50386 176700 79455
rect 176764 51066 176792 79494
rect 176856 78305 176884 79614
rect 176842 78296 176898 78305
rect 176842 78231 176898 78240
rect 176844 75132 176896 75138
rect 176844 75074 176896 75080
rect 176856 61946 176884 75074
rect 176948 68882 176976 79716
rect 177040 74934 177068 79784
rect 177178 79676 177206 80036
rect 177270 79812 177298 80036
rect 177362 79971 177390 80036
rect 177348 79962 177404 79971
rect 177348 79897 177404 79906
rect 177454 79812 177482 80036
rect 177546 79971 177574 80036
rect 177532 79962 177588 79971
rect 177532 79897 177588 79906
rect 177638 79914 177666 80036
rect 177638 79886 177712 79914
rect 177580 79824 177632 79830
rect 177270 79784 177344 79812
rect 177454 79801 177528 79812
rect 177454 79792 177542 79801
rect 177454 79784 177486 79792
rect 177316 79778 177344 79784
rect 177316 79750 177390 79778
rect 177362 79744 177390 79750
rect 177362 79716 177436 79744
rect 177580 79766 177632 79772
rect 177486 79727 177542 79736
rect 177132 79648 177206 79676
rect 177132 75138 177160 79648
rect 177408 77994 177436 79716
rect 177488 79620 177540 79626
rect 177488 79562 177540 79568
rect 177396 77988 177448 77994
rect 177396 77930 177448 77936
rect 177212 77920 177264 77926
rect 177210 77888 177212 77897
rect 177264 77888 177266 77897
rect 177210 77823 177266 77832
rect 177304 77376 177356 77382
rect 177304 77318 177356 77324
rect 177120 75132 177172 75138
rect 177120 75074 177172 75080
rect 177028 74928 177080 74934
rect 177028 74870 177080 74876
rect 176936 68876 176988 68882
rect 176936 68818 176988 68824
rect 176844 61940 176896 61946
rect 176844 61882 176896 61888
rect 176752 51060 176804 51066
rect 176752 51002 176804 51008
rect 176660 50380 176712 50386
rect 176660 50322 176712 50328
rect 177316 29714 177344 77318
rect 177500 77314 177528 79562
rect 177592 79257 177620 79766
rect 177684 79529 177712 79886
rect 177670 79520 177726 79529
rect 177670 79455 177726 79464
rect 177578 79248 177634 79257
rect 177578 79183 177634 79192
rect 177488 77308 177540 77314
rect 177488 77250 177540 77256
rect 177488 74928 177540 74934
rect 177488 74870 177540 74876
rect 177500 46918 177528 74870
rect 177684 47598 177712 79455
rect 177776 79354 177804 80038
rect 177856 80028 177908 80034
rect 177908 79988 177988 80016
rect 177856 79970 177908 79976
rect 177856 79892 177908 79898
rect 177856 79834 177908 79840
rect 177764 79348 177816 79354
rect 177764 79290 177816 79296
rect 177868 78418 177896 79834
rect 177776 78390 177896 78418
rect 177776 75138 177804 78390
rect 177854 78296 177910 78305
rect 177854 78231 177910 78240
rect 177868 77994 177896 78231
rect 177856 77988 177908 77994
rect 177856 77930 177908 77936
rect 177764 75132 177816 75138
rect 177764 75074 177816 75080
rect 177672 47592 177724 47598
rect 177672 47534 177724 47540
rect 177488 46912 177540 46918
rect 177488 46854 177540 46860
rect 177776 35222 177804 75074
rect 177764 35216 177816 35222
rect 177764 35158 177816 35164
rect 177868 33794 177896 77930
rect 177960 77042 177988 79988
rect 178052 79490 178080 80310
rect 178144 79694 178172 80407
rect 178500 80164 178552 80170
rect 178500 80106 178552 80112
rect 178224 79756 178276 79762
rect 178224 79698 178276 79704
rect 178132 79688 178184 79694
rect 178132 79630 178184 79636
rect 178040 79484 178092 79490
rect 178040 79426 178092 79432
rect 178236 78810 178264 79698
rect 178224 78804 178276 78810
rect 178224 78746 178276 78752
rect 178038 77616 178094 77625
rect 178038 77551 178094 77560
rect 177948 77036 178000 77042
rect 177948 76978 178000 76984
rect 177856 33788 177908 33794
rect 177856 33730 177908 33736
rect 177304 29708 177356 29714
rect 177304 29650 177356 29656
rect 177960 18630 177988 76978
rect 178052 75206 178080 77551
rect 178512 75750 178540 80106
rect 178592 80028 178644 80034
rect 178592 79970 178644 79976
rect 178604 76945 178632 79970
rect 178788 79558 178816 80582
rect 179340 80238 179368 80679
rect 179616 80442 179644 80679
rect 179604 80436 179656 80442
rect 179604 80378 179656 80384
rect 179892 80306 179920 80679
rect 181442 80472 181498 80481
rect 181442 80407 181498 80416
rect 179880 80300 179932 80306
rect 179880 80242 179932 80248
rect 179328 80232 179380 80238
rect 181456 80209 181484 80407
rect 179328 80174 179380 80180
rect 181442 80200 181498 80209
rect 181442 80135 181498 80144
rect 181168 80096 181220 80102
rect 179326 80064 179382 80073
rect 181168 80038 181220 80044
rect 179326 79999 179382 80008
rect 178776 79552 178828 79558
rect 178776 79494 178828 79500
rect 178960 78056 179012 78062
rect 178960 77998 179012 78004
rect 178776 77852 178828 77858
rect 178776 77794 178828 77800
rect 178590 76936 178646 76945
rect 178590 76871 178646 76880
rect 178684 76492 178736 76498
rect 178684 76434 178736 76440
rect 178500 75744 178552 75750
rect 178500 75686 178552 75692
rect 178040 75200 178092 75206
rect 178040 75142 178092 75148
rect 178038 72448 178094 72457
rect 178038 72383 178094 72392
rect 177948 18624 178000 18630
rect 177948 18566 178000 18572
rect 178052 16574 178080 72383
rect 178052 16546 178632 16574
rect 176568 6248 176620 6254
rect 176568 6190 176620 6196
rect 175832 6180 175884 6186
rect 175832 6122 175884 6128
rect 173900 4820 173952 4826
rect 173900 4762 173952 4768
rect 173256 3596 173308 3602
rect 173256 3538 173308 3544
rect 177856 3596 177908 3602
rect 177856 3538 177908 3544
rect 175464 3528 175516 3534
rect 175464 3470 175516 3476
rect 174268 3188 174320 3194
rect 174268 3130 174320 3136
rect 174280 480 174308 3130
rect 175476 480 175504 3470
rect 176660 3460 176712 3466
rect 176660 3402 176712 3408
rect 176672 480 176700 3402
rect 177868 480 177896 3538
rect 164854 354 164966 480
rect 164528 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3466 178724 76434
rect 178788 13258 178816 77794
rect 178868 77512 178920 77518
rect 178868 77454 178920 77460
rect 178880 27062 178908 77454
rect 178972 33114 179000 77998
rect 179234 77888 179290 77897
rect 179234 77823 179290 77832
rect 179248 70394 179276 77823
rect 179340 77382 179368 79999
rect 181074 79520 181130 79529
rect 181074 79455 181130 79464
rect 179510 78976 179566 78985
rect 179510 78911 179566 78920
rect 180890 78976 180946 78985
rect 181088 78946 181116 79455
rect 181180 78985 181208 80038
rect 182086 79792 182142 79801
rect 182086 79727 182142 79736
rect 181166 78976 181222 78985
rect 180890 78911 180946 78920
rect 181076 78940 181128 78946
rect 179524 78742 179552 78911
rect 180904 78878 180932 78911
rect 181166 78911 181222 78920
rect 181076 78882 181128 78888
rect 180892 78872 180944 78878
rect 180892 78814 180944 78820
rect 179512 78736 179564 78742
rect 179512 78678 179564 78684
rect 179328 77376 179380 77382
rect 179328 77318 179380 77324
rect 179326 77208 179382 77217
rect 179326 77143 179382 77152
rect 179340 76974 179368 77143
rect 179328 76968 179380 76974
rect 179328 76910 179380 76916
rect 179340 75954 179368 76910
rect 179328 75948 179380 75954
rect 179328 75890 179380 75896
rect 179524 71126 179552 78678
rect 180800 78056 180852 78062
rect 180800 77998 180852 78004
rect 180812 77586 180840 77998
rect 180800 77580 180852 77586
rect 180800 77522 180852 77528
rect 180062 77208 180118 77217
rect 180062 77143 180118 77152
rect 180076 76022 180104 77143
rect 180064 76016 180116 76022
rect 180064 75958 180116 75964
rect 180064 75064 180116 75070
rect 180064 75006 180116 75012
rect 179420 71120 179472 71126
rect 179420 71062 179472 71068
rect 179512 71120 179564 71126
rect 179512 71062 179564 71068
rect 179248 70366 179368 70394
rect 178960 33108 179012 33114
rect 178960 33050 179012 33056
rect 178868 27056 178920 27062
rect 178868 26998 178920 27004
rect 179340 14618 179368 70366
rect 179432 16574 179460 71062
rect 179432 16546 180012 16574
rect 179328 14612 179380 14618
rect 179328 14554 179380 14560
rect 178776 13252 178828 13258
rect 178776 13194 178828 13200
rect 179984 3482 180012 16546
rect 180076 3602 180104 75006
rect 180800 74996 180852 75002
rect 180800 74938 180852 74944
rect 180812 16574 180840 74938
rect 180904 70990 180932 78814
rect 181444 78600 181496 78606
rect 181444 78542 181496 78548
rect 181456 77450 181484 78542
rect 181536 77920 181588 77926
rect 181534 77888 181536 77897
rect 181588 77888 181590 77897
rect 181534 77823 181590 77832
rect 182100 77489 182128 79727
rect 186320 78872 186372 78878
rect 186320 78814 186372 78820
rect 186332 78538 186360 78814
rect 186412 78804 186464 78810
rect 186412 78746 186464 78752
rect 186320 78532 186372 78538
rect 186320 78474 186372 78480
rect 186424 78470 186452 78746
rect 186412 78464 186464 78470
rect 186412 78406 186464 78412
rect 183100 78396 183152 78402
rect 183100 78338 183152 78344
rect 182086 77480 182142 77489
rect 181444 77444 181496 77450
rect 182086 77415 182142 77424
rect 181444 77386 181496 77392
rect 181444 76628 181496 76634
rect 181444 76570 181496 76576
rect 180892 70984 180944 70990
rect 180892 70926 180944 70932
rect 180812 16546 181024 16574
rect 180064 3596 180116 3602
rect 180064 3538 180116 3544
rect 178684 3460 178736 3466
rect 179984 3454 180288 3482
rect 178684 3402 178736 3408
rect 180260 480 180288 3454
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 181456 3738 181484 76570
rect 182824 75676 182876 75682
rect 182824 75618 182876 75624
rect 181536 69692 181588 69698
rect 181536 69634 181588 69640
rect 181444 3732 181496 3738
rect 181444 3674 181496 3680
rect 181548 3602 181576 69634
rect 181536 3596 181588 3602
rect 181536 3538 181588 3544
rect 182548 3596 182600 3602
rect 182548 3538 182600 3544
rect 182560 480 182588 3538
rect 182836 3126 182864 75618
rect 182914 70000 182970 70009
rect 182914 69935 182970 69944
rect 182824 3120 182876 3126
rect 182824 3062 182876 3068
rect 182928 3058 182956 69935
rect 183006 68912 183062 68921
rect 183006 68847 183062 68856
rect 183020 68814 183048 68847
rect 183008 68808 183060 68814
rect 183008 68750 183060 68756
rect 183008 64184 183060 64190
rect 183008 64126 183060 64132
rect 183020 3602 183048 64126
rect 183112 31142 183140 78338
rect 183652 78124 183704 78130
rect 183652 78066 183704 78072
rect 183560 75744 183612 75750
rect 183560 75686 183612 75692
rect 183572 75041 183600 75686
rect 183558 75032 183614 75041
rect 183558 74967 183614 74976
rect 183664 71738 183692 78066
rect 185582 77480 185638 77489
rect 185582 77415 185638 77424
rect 183652 71732 183704 71738
rect 183652 71674 183704 71680
rect 185032 71120 185084 71126
rect 185032 71062 185084 71068
rect 183468 68808 183520 68814
rect 183468 68750 183520 68756
rect 183480 67726 183508 68750
rect 184202 68368 184258 68377
rect 184202 68303 184258 68312
rect 183468 67720 183520 67726
rect 183468 67662 183520 67668
rect 183560 65544 183612 65550
rect 183560 65486 183612 65492
rect 183100 31136 183152 31142
rect 183100 31078 183152 31084
rect 183572 16574 183600 65486
rect 183572 16546 183784 16574
rect 183008 3596 183060 3602
rect 183008 3538 183060 3544
rect 182916 3052 182968 3058
rect 182916 2994 182968 3000
rect 183756 480 183784 16546
rect 184216 3806 184244 68303
rect 185044 6914 185072 71062
rect 185596 8974 185624 77415
rect 186320 60036 186372 60042
rect 186320 59978 186372 59984
rect 186332 16574 186360 59978
rect 186608 57905 186636 195230
rect 186700 76537 186728 197882
rect 186792 81054 186820 200126
rect 187516 198892 187568 198898
rect 187516 198834 187568 198840
rect 187056 198620 187108 198626
rect 187056 198562 187108 198568
rect 186872 198552 186924 198558
rect 186872 198494 186924 198500
rect 186780 81048 186832 81054
rect 186780 80990 186832 80996
rect 186792 80850 186820 80990
rect 186780 80844 186832 80850
rect 186780 80786 186832 80792
rect 186884 80209 186912 198494
rect 186964 198348 187016 198354
rect 186964 198290 187016 198296
rect 186870 80200 186926 80209
rect 186870 80135 186926 80144
rect 186976 78878 187004 198290
rect 186964 78872 187016 78878
rect 186964 78814 187016 78820
rect 187068 78810 187096 198562
rect 187424 197872 187476 197878
rect 187424 197814 187476 197820
rect 187148 149048 187200 149054
rect 187148 148990 187200 148996
rect 187056 78804 187108 78810
rect 187056 78746 187108 78752
rect 186686 76528 186742 76537
rect 186686 76463 186742 76472
rect 186700 68338 186728 76463
rect 187160 71194 187188 148990
rect 187240 141976 187292 141982
rect 187240 141918 187292 141924
rect 187252 72282 187280 141918
rect 187330 139224 187386 139233
rect 187330 139159 187386 139168
rect 187344 75857 187372 139159
rect 187436 138145 187464 197814
rect 187528 138281 187556 198834
rect 187712 142594 187740 273226
rect 188252 262676 188304 262682
rect 188252 262618 188304 262624
rect 187884 200388 187936 200394
rect 187884 200330 187936 200336
rect 187792 198960 187844 198966
rect 187792 198902 187844 198908
rect 187700 142588 187752 142594
rect 187700 142530 187752 142536
rect 187514 138272 187570 138281
rect 187514 138207 187570 138216
rect 187422 138136 187478 138145
rect 187422 138071 187478 138080
rect 187424 81252 187476 81258
rect 187424 81194 187476 81200
rect 187436 80918 187464 81194
rect 187516 81116 187568 81122
rect 187516 81058 187568 81064
rect 187424 80912 187476 80918
rect 187424 80854 187476 80860
rect 187422 80200 187478 80209
rect 187422 80135 187478 80144
rect 187330 75848 187386 75857
rect 187330 75783 187386 75792
rect 187240 72276 187292 72282
rect 187240 72218 187292 72224
rect 187148 71188 187200 71194
rect 187148 71130 187200 71136
rect 187436 69737 187464 80135
rect 187528 77722 187556 81058
rect 187700 78736 187752 78742
rect 187700 78678 187752 78684
rect 187516 77716 187568 77722
rect 187516 77658 187568 77664
rect 187712 77489 187740 78678
rect 187698 77480 187754 77489
rect 187698 77415 187754 77424
rect 187700 75608 187752 75614
rect 187700 75550 187752 75556
rect 187422 69728 187478 69737
rect 187422 69663 187478 69672
rect 186688 68332 186740 68338
rect 186688 68274 186740 68280
rect 186962 62112 187018 62121
rect 186962 62047 187018 62056
rect 186976 61878 187004 62047
rect 186964 61872 187016 61878
rect 186964 61814 187016 61820
rect 186976 60858 187004 61814
rect 186964 60852 187016 60858
rect 186964 60794 187016 60800
rect 186594 57896 186650 57905
rect 186594 57831 186650 57840
rect 187712 16574 187740 75550
rect 187804 63209 187832 198902
rect 187896 66201 187924 200330
rect 188160 199572 188212 199578
rect 188160 199514 188212 199520
rect 187976 198416 188028 198422
rect 187976 198358 188028 198364
rect 187988 75818 188016 198358
rect 188068 198280 188120 198286
rect 188068 198222 188120 198228
rect 187976 75812 188028 75818
rect 187976 75754 188028 75760
rect 188080 75177 188108 198222
rect 188172 80782 188200 199514
rect 188264 144362 188292 262618
rect 188988 260432 189040 260438
rect 188988 260374 189040 260380
rect 189000 259418 189028 260374
rect 188988 259412 189040 259418
rect 188988 259354 189040 259360
rect 189092 200705 189120 282882
rect 190460 265600 190512 265606
rect 190460 265542 190512 265548
rect 189172 262268 189224 262274
rect 189172 262210 189224 262216
rect 189078 200696 189134 200705
rect 189078 200631 189134 200640
rect 189080 199164 189132 199170
rect 189080 199106 189132 199112
rect 188344 198688 188396 198694
rect 188344 198630 188396 198636
rect 188252 144356 188304 144362
rect 188252 144298 188304 144304
rect 188250 139360 188306 139369
rect 188250 139295 188306 139304
rect 188160 80776 188212 80782
rect 188160 80718 188212 80724
rect 188066 75168 188122 75177
rect 188066 75103 188122 75112
rect 187882 66192 187938 66201
rect 187882 66127 187938 66136
rect 187896 65929 187924 66127
rect 187882 65920 187938 65929
rect 187882 65855 187938 65864
rect 187790 63200 187846 63209
rect 187790 63135 187846 63144
rect 188264 59129 188292 139295
rect 188356 78742 188384 198630
rect 188436 198212 188488 198218
rect 188436 198154 188488 198160
rect 188448 80481 188476 198154
rect 188528 178084 188580 178090
rect 188528 178026 188580 178032
rect 188540 144294 188568 178026
rect 188528 144288 188580 144294
rect 188528 144230 188580 144236
rect 188620 139596 188672 139602
rect 188620 139538 188672 139544
rect 188526 127664 188582 127673
rect 188526 127599 188582 127608
rect 188434 80472 188490 80481
rect 188434 80407 188490 80416
rect 188344 78736 188396 78742
rect 188344 78678 188396 78684
rect 188448 71369 188476 80407
rect 188434 71360 188490 71369
rect 188434 71295 188490 71304
rect 188344 71120 188396 71126
rect 188344 71062 188396 71068
rect 188356 70990 188384 71062
rect 188344 70984 188396 70990
rect 188344 70926 188396 70932
rect 188540 69766 188568 127599
rect 188632 74458 188660 139538
rect 188620 74452 188672 74458
rect 188620 74394 188672 74400
rect 188528 69760 188580 69766
rect 188528 69702 188580 69708
rect 189092 63073 189120 199106
rect 189184 198830 189212 262210
rect 189724 261588 189776 261594
rect 189724 261530 189776 261536
rect 189632 260092 189684 260098
rect 189632 260034 189684 260040
rect 189540 260024 189592 260030
rect 189540 259966 189592 259972
rect 189356 259888 189408 259894
rect 189356 259830 189408 259836
rect 189172 198824 189224 198830
rect 189172 198766 189224 198772
rect 189264 195220 189316 195226
rect 189264 195162 189316 195168
rect 189172 195016 189224 195022
rect 189172 194958 189224 194964
rect 189184 70786 189212 194958
rect 189172 70780 189224 70786
rect 189172 70722 189224 70728
rect 189276 70666 189304 195162
rect 189368 141438 189396 259830
rect 189446 259584 189502 259593
rect 189446 259519 189502 259528
rect 189460 142118 189488 259519
rect 189552 143313 189580 259966
rect 189538 143304 189594 143313
rect 189538 143239 189594 143248
rect 189644 142798 189672 260034
rect 189736 193186 189764 261530
rect 190472 200802 190500 265542
rect 190828 265532 190880 265538
rect 190828 265474 190880 265480
rect 190552 262404 190604 262410
rect 190552 262346 190604 262352
rect 190460 200796 190512 200802
rect 190460 200738 190512 200744
rect 190564 199510 190592 262346
rect 190644 262336 190696 262342
rect 190644 262278 190696 262284
rect 190552 199504 190604 199510
rect 190552 199446 190604 199452
rect 190656 199442 190684 262278
rect 190736 200252 190788 200258
rect 190736 200194 190788 200200
rect 190644 199436 190696 199442
rect 190644 199378 190696 199384
rect 189816 199232 189868 199238
rect 189816 199174 189868 199180
rect 189724 193180 189776 193186
rect 189724 193122 189776 193128
rect 189724 165640 189776 165646
rect 189724 165582 189776 165588
rect 189736 144226 189764 165582
rect 189724 144220 189776 144226
rect 189724 144162 189776 144168
rect 189632 142792 189684 142798
rect 189632 142734 189684 142740
rect 189448 142112 189500 142118
rect 189448 142054 189500 142060
rect 189356 141432 189408 141438
rect 189356 141374 189408 141380
rect 189724 140412 189776 140418
rect 189724 140354 189776 140360
rect 189540 140344 189592 140350
rect 189540 140286 189592 140292
rect 189552 76702 189580 140286
rect 189632 139936 189684 139942
rect 189632 139878 189684 139884
rect 189644 77110 189672 139878
rect 189632 77104 189684 77110
rect 189632 77046 189684 77052
rect 189644 76702 189672 77046
rect 189540 76696 189592 76702
rect 189540 76638 189592 76644
rect 189632 76696 189684 76702
rect 189632 76638 189684 76644
rect 189736 76362 189764 140354
rect 189828 139777 189856 199174
rect 190644 195968 190696 195974
rect 190644 195910 190696 195916
rect 190460 195492 190512 195498
rect 190460 195434 190512 195440
rect 190000 145648 190052 145654
rect 190000 145590 190052 145596
rect 189908 140004 189960 140010
rect 189908 139946 189960 139952
rect 189814 139768 189870 139777
rect 189814 139703 189870 139712
rect 189816 139460 189868 139466
rect 189816 139402 189868 139408
rect 189828 79694 189856 139402
rect 189816 79688 189868 79694
rect 189816 79630 189868 79636
rect 189920 79354 189948 139946
rect 189908 79348 189960 79354
rect 189908 79290 189960 79296
rect 189724 76356 189776 76362
rect 189724 76298 189776 76304
rect 190012 72418 190040 145590
rect 190092 143336 190144 143342
rect 190092 143278 190144 143284
rect 190184 143336 190236 143342
rect 190184 143278 190236 143284
rect 190104 73030 190132 143278
rect 190196 143070 190224 143278
rect 190184 143064 190236 143070
rect 190184 143006 190236 143012
rect 190092 73024 190144 73030
rect 190092 72966 190144 72972
rect 190000 72412 190052 72418
rect 190000 72354 190052 72360
rect 189356 70780 189408 70786
rect 189356 70722 189408 70728
rect 189184 70638 189304 70666
rect 189184 68950 189212 70638
rect 189172 68944 189224 68950
rect 189172 68886 189224 68892
rect 189184 68406 189212 68886
rect 189172 68400 189224 68406
rect 189172 68342 189224 68348
rect 189170 67552 189226 67561
rect 189170 67487 189226 67496
rect 189184 66298 189212 67487
rect 189368 67425 189396 70722
rect 189722 68232 189778 68241
rect 189722 68167 189778 68176
rect 189354 67416 189410 67425
rect 189354 67351 189410 67360
rect 189172 66292 189224 66298
rect 189172 66234 189224 66240
rect 189078 63064 189134 63073
rect 189078 62999 189134 63008
rect 188250 59120 188306 59129
rect 188250 59055 188306 59064
rect 189736 16574 189764 68167
rect 189906 67416 189962 67425
rect 189906 67351 189962 67360
rect 189920 67017 189948 67351
rect 189906 67008 189962 67017
rect 189906 66943 189962 66952
rect 190472 50833 190500 195434
rect 190552 195356 190604 195362
rect 190552 195298 190604 195304
rect 190564 57633 190592 195298
rect 190656 61985 190684 195910
rect 190748 79626 190776 200194
rect 190840 144838 190868 265474
rect 194876 265464 194928 265470
rect 194876 265406 194928 265412
rect 192024 265328 192076 265334
rect 192024 265270 192076 265276
rect 190920 263628 190972 263634
rect 190920 263570 190972 263576
rect 190828 144832 190880 144838
rect 190828 144774 190880 144780
rect 190932 143041 190960 263570
rect 191012 263492 191064 263498
rect 191012 263434 191064 263440
rect 191024 262614 191052 263434
rect 191840 263424 191892 263430
rect 191840 263366 191892 263372
rect 191012 262608 191064 262614
rect 191012 262550 191064 262556
rect 191024 262313 191052 262550
rect 191852 262546 191880 263366
rect 191840 262540 191892 262546
rect 191840 262482 191892 262488
rect 191852 262313 191880 262482
rect 191010 262304 191066 262313
rect 191010 262239 191066 262248
rect 191838 262304 191894 262313
rect 191838 262239 191894 262248
rect 191196 260228 191248 260234
rect 191196 260170 191248 260176
rect 191012 259956 191064 259962
rect 191012 259898 191064 259904
rect 190918 143032 190974 143041
rect 190918 142967 190974 142976
rect 191024 142934 191052 259898
rect 191104 259752 191156 259758
rect 191104 259694 191156 259700
rect 191012 142928 191064 142934
rect 191012 142870 191064 142876
rect 191116 142866 191144 259694
rect 191208 143138 191236 260170
rect 191378 259992 191434 260001
rect 191378 259927 191434 259936
rect 191288 144152 191340 144158
rect 191288 144094 191340 144100
rect 191196 143132 191248 143138
rect 191196 143074 191248 143080
rect 191104 142860 191156 142866
rect 191104 142802 191156 142808
rect 190920 141160 190972 141166
rect 190920 141102 190972 141108
rect 190828 140752 190880 140758
rect 190826 140720 190828 140729
rect 190880 140720 190882 140729
rect 190826 140655 190882 140664
rect 190826 138680 190882 138689
rect 190826 138615 190882 138624
rect 190736 79620 190788 79626
rect 190736 79562 190788 79568
rect 190642 61976 190698 61985
rect 190642 61911 190698 61920
rect 190550 57624 190606 57633
rect 190550 57559 190606 57568
rect 190840 56409 190868 138615
rect 190932 66230 190960 141102
rect 191196 140956 191248 140962
rect 191196 140898 191248 140904
rect 191102 138544 191158 138553
rect 191102 138479 191158 138488
rect 191116 72486 191144 138479
rect 191208 77178 191236 140898
rect 191300 79762 191328 144094
rect 191392 143177 191420 259927
rect 191932 196512 191984 196518
rect 191932 196454 191984 196460
rect 191840 196444 191892 196450
rect 191840 196386 191892 196392
rect 191472 143472 191524 143478
rect 191472 143414 191524 143420
rect 191378 143168 191434 143177
rect 191378 143103 191434 143112
rect 191288 79756 191340 79762
rect 191288 79698 191340 79704
rect 191196 77172 191248 77178
rect 191196 77114 191248 77120
rect 191484 74497 191512 143414
rect 191748 77172 191800 77178
rect 191748 77114 191800 77120
rect 191760 76634 191788 77114
rect 191748 76628 191800 76634
rect 191748 76570 191800 76576
rect 191470 74488 191526 74497
rect 191470 74423 191526 74432
rect 191484 73817 191512 74423
rect 191470 73808 191526 73817
rect 191470 73743 191526 73752
rect 191104 72480 191156 72486
rect 191104 72422 191156 72428
rect 190920 66224 190972 66230
rect 190920 66166 190972 66172
rect 191748 66224 191800 66230
rect 191748 66166 191800 66172
rect 191760 65550 191788 66166
rect 191748 65544 191800 65550
rect 191748 65486 191800 65492
rect 191746 61976 191802 61985
rect 191746 61911 191802 61920
rect 191760 61577 191788 61911
rect 191746 61568 191802 61577
rect 191746 61503 191802 61512
rect 190826 56400 190882 56409
rect 190826 56335 190882 56344
rect 191852 55049 191880 196386
rect 191944 58857 191972 196454
rect 192036 141642 192064 265270
rect 193404 264988 193456 264994
rect 193404 264930 193456 264936
rect 192484 263152 192536 263158
rect 192484 263094 192536 263100
rect 192300 263016 192352 263022
rect 192300 262958 192352 262964
rect 192208 262812 192260 262818
rect 192208 262754 192260 262760
rect 192116 200320 192168 200326
rect 192116 200262 192168 200268
rect 192024 141636 192076 141642
rect 192024 141578 192076 141584
rect 192128 84194 192156 200262
rect 192220 141506 192248 262754
rect 192312 141574 192340 262958
rect 192392 260296 192444 260302
rect 192392 260238 192444 260244
rect 192404 143206 192432 260238
rect 192496 145450 192524 263094
rect 193220 199028 193272 199034
rect 193220 198970 193272 198976
rect 192760 147416 192812 147422
rect 192760 147358 192812 147364
rect 192484 145444 192536 145450
rect 192484 145386 192536 145392
rect 192392 143200 192444 143206
rect 192392 143142 192444 143148
rect 192300 141568 192352 141574
rect 192300 141510 192352 141516
rect 192208 141500 192260 141506
rect 192208 141442 192260 141448
rect 192392 140276 192444 140282
rect 192392 140218 192444 140224
rect 192298 138408 192354 138417
rect 192298 138343 192354 138352
rect 192036 84166 192156 84194
rect 192036 79082 192064 84166
rect 192024 79076 192076 79082
rect 192024 79018 192076 79024
rect 192312 71262 192340 138343
rect 192404 73778 192432 140218
rect 192576 140208 192628 140214
rect 192576 140150 192628 140156
rect 192588 76906 192616 140150
rect 192668 139868 192720 139874
rect 192668 139810 192720 139816
rect 192680 81122 192708 139810
rect 192668 81116 192720 81122
rect 192668 81058 192720 81064
rect 192576 76900 192628 76906
rect 192576 76842 192628 76848
rect 192772 76838 192800 147358
rect 192852 146872 192904 146878
rect 192852 146814 192904 146820
rect 192864 78606 192892 146814
rect 192944 145784 192996 145790
rect 192944 145726 192996 145732
rect 192956 79150 192984 145726
rect 192944 79144 192996 79150
rect 192944 79086 192996 79092
rect 192852 78600 192904 78606
rect 192852 78542 192904 78548
rect 192760 76832 192812 76838
rect 192760 76774 192812 76780
rect 192392 73772 192444 73778
rect 192392 73714 192444 73720
rect 192300 71256 192352 71262
rect 192300 71198 192352 71204
rect 193232 63510 193260 198970
rect 193312 195900 193364 195906
rect 193312 195842 193364 195848
rect 193220 63504 193272 63510
rect 193220 63446 193272 63452
rect 193232 62898 193260 63446
rect 193220 62892 193272 62898
rect 193220 62834 193272 62840
rect 193324 60722 193352 195842
rect 193416 145722 193444 264930
rect 193588 262744 193640 262750
rect 193588 262686 193640 262692
rect 193496 260500 193548 260506
rect 193496 260442 193548 260448
rect 193404 145716 193456 145722
rect 193404 145658 193456 145664
rect 193402 144936 193458 144945
rect 193402 144871 193458 144880
rect 193416 144498 193444 144871
rect 193404 144492 193456 144498
rect 193404 144434 193456 144440
rect 193508 141710 193536 260442
rect 193600 144634 193628 262686
rect 193772 261316 193824 261322
rect 193772 261258 193824 261264
rect 193680 261112 193732 261118
rect 193680 261054 193732 261060
rect 193588 144628 193640 144634
rect 193588 144570 193640 144576
rect 193692 144430 193720 261054
rect 193784 156670 193812 261258
rect 194692 197260 194744 197266
rect 194692 197202 194744 197208
rect 194600 196852 194652 196858
rect 194600 196794 194652 196800
rect 193864 192976 193916 192982
rect 193864 192918 193916 192924
rect 193772 156664 193824 156670
rect 193772 156606 193824 156612
rect 193680 144424 193732 144430
rect 193680 144366 193732 144372
rect 193772 141908 193824 141914
rect 193772 141850 193824 141856
rect 193496 141704 193548 141710
rect 193496 141646 193548 141652
rect 193588 140548 193640 140554
rect 193588 140490 193640 140496
rect 193402 138952 193458 138961
rect 193402 138887 193458 138896
rect 193312 60716 193364 60722
rect 193312 60658 193364 60664
rect 191930 58848 191986 58857
rect 191930 58783 191986 58792
rect 193312 58744 193364 58750
rect 193312 58686 193364 58692
rect 191838 55040 191894 55049
rect 191838 54975 191894 54984
rect 191852 54777 191880 54975
rect 191838 54768 191894 54777
rect 191838 54703 191894 54712
rect 191840 51740 191892 51746
rect 191840 51682 191892 51688
rect 190458 50824 190514 50833
rect 190458 50759 190514 50768
rect 191852 16574 191880 51682
rect 193324 16574 193352 58686
rect 193416 54913 193444 138887
rect 193600 66065 193628 140490
rect 193586 66056 193642 66065
rect 193586 65991 193642 66000
rect 193784 57497 193812 141850
rect 193876 79286 193904 192918
rect 193956 156664 194008 156670
rect 193956 156606 194008 156612
rect 193968 146130 193996 156606
rect 194140 148300 194192 148306
rect 194140 148242 194192 148248
rect 194048 147280 194100 147286
rect 194048 147222 194100 147228
rect 193956 146124 194008 146130
rect 193956 146066 194008 146072
rect 193956 140616 194008 140622
rect 193956 140558 194008 140564
rect 193864 79280 193916 79286
rect 193864 79222 193916 79228
rect 193968 70922 193996 140558
rect 194060 79490 194088 147222
rect 194048 79484 194100 79490
rect 194048 79426 194100 79432
rect 194152 77926 194180 148242
rect 194232 144560 194284 144566
rect 194232 144502 194284 144508
rect 194140 77920 194192 77926
rect 194140 77862 194192 77868
rect 194244 71398 194272 144502
rect 194232 71392 194284 71398
rect 194232 71334 194284 71340
rect 193956 70916 194008 70922
rect 193956 70858 194008 70864
rect 193862 66872 193918 66881
rect 193862 66807 193918 66816
rect 193770 57488 193826 57497
rect 193770 57423 193826 57432
rect 193402 54904 193458 54913
rect 193402 54839 193458 54848
rect 193416 54641 193444 54839
rect 193402 54632 193458 54641
rect 193402 54567 193458 54576
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 189736 16546 189856 16574
rect 191852 16546 192064 16574
rect 193324 16546 193812 16574
rect 185584 8968 185636 8974
rect 185584 8910 185636 8916
rect 185044 6886 186176 6914
rect 184204 3800 184256 3806
rect 184204 3742 184256 3748
rect 184940 3120 184992 3126
rect 184940 3062 184992 3068
rect 184952 480 184980 3062
rect 186148 480 186176 6886
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 189828 3670 189856 16546
rect 189816 3664 189868 3670
rect 189816 3606 189868 3612
rect 190828 3596 190880 3602
rect 190828 3538 190880 3544
rect 189724 3052 189776 3058
rect 189724 2994 189776 3000
rect 189736 480 189764 2994
rect 190840 480 190868 3538
rect 192036 480 192064 16546
rect 193220 3664 193272 3670
rect 193220 3606 193272 3612
rect 193232 480 193260 3606
rect 193784 3482 193812 16546
rect 193876 3602 193904 66807
rect 194506 66056 194562 66065
rect 194506 65991 194562 66000
rect 194520 65793 194548 65991
rect 194506 65784 194562 65793
rect 194506 65719 194562 65728
rect 194508 60716 194560 60722
rect 194508 60658 194560 60664
rect 194520 60042 194548 60658
rect 194508 60036 194560 60042
rect 194508 59978 194560 59984
rect 194612 47705 194640 196794
rect 194704 52329 194732 197202
rect 194784 197192 194836 197198
rect 194784 197134 194836 197140
rect 194796 53689 194824 197134
rect 194888 145518 194916 265406
rect 196440 265396 196492 265402
rect 196440 265338 196492 265344
rect 196256 265124 196308 265130
rect 196256 265066 196308 265072
rect 194968 263696 195020 263702
rect 194968 263638 195020 263644
rect 194876 145512 194928 145518
rect 194876 145454 194928 145460
rect 194980 144770 195008 263638
rect 195060 260976 195112 260982
rect 195060 260918 195112 260924
rect 195072 146266 195100 260918
rect 195244 259616 195296 259622
rect 195244 259558 195296 259564
rect 195152 195628 195204 195634
rect 195152 195570 195204 195576
rect 195060 146260 195112 146266
rect 195060 146202 195112 146208
rect 195060 145920 195112 145926
rect 195060 145862 195112 145868
rect 194968 144764 195020 144770
rect 194968 144706 195020 144712
rect 194966 139088 195022 139097
rect 194966 139023 195022 139032
rect 194980 71670 195008 139023
rect 195072 79121 195100 145862
rect 195164 80714 195192 195570
rect 195256 146062 195284 259558
rect 195336 198144 195388 198150
rect 195336 198086 195388 198092
rect 195348 146985 195376 198086
rect 196072 196988 196124 196994
rect 196072 196930 196124 196936
rect 195980 195424 196032 195430
rect 195980 195366 196032 195372
rect 195428 148980 195480 148986
rect 195428 148922 195480 148928
rect 195334 146976 195390 146985
rect 195334 146911 195390 146920
rect 195244 146056 195296 146062
rect 195244 145998 195296 146004
rect 195336 145988 195388 145994
rect 195336 145930 195388 145936
rect 195348 81297 195376 145930
rect 195334 81288 195390 81297
rect 195334 81223 195390 81232
rect 195152 80708 195204 80714
rect 195152 80650 195204 80656
rect 195058 79112 195114 79121
rect 195058 79047 195114 79056
rect 194968 71664 195020 71670
rect 194968 71606 195020 71612
rect 195440 71330 195468 148922
rect 195520 147144 195572 147150
rect 195520 147086 195572 147092
rect 195532 81161 195560 147086
rect 195518 81152 195574 81161
rect 195518 81087 195574 81096
rect 195428 71324 195480 71330
rect 195428 71266 195480 71272
rect 194782 53680 194838 53689
rect 194782 53615 194838 53624
rect 194796 53281 194824 53615
rect 194782 53272 194838 53281
rect 194782 53207 194838 53216
rect 194690 52320 194746 52329
rect 194690 52255 194746 52264
rect 194704 51921 194732 52255
rect 194690 51912 194746 51921
rect 194690 51847 194746 51856
rect 195992 49473 196020 195366
rect 196084 64874 196112 196930
rect 196164 196648 196216 196654
rect 196164 196590 196216 196596
rect 196176 66745 196204 196590
rect 196268 144702 196296 265066
rect 196348 262472 196400 262478
rect 196348 262414 196400 262420
rect 196256 144696 196308 144702
rect 196256 144638 196308 144644
rect 196360 141846 196388 262414
rect 196452 147626 196480 265338
rect 197636 265260 197688 265266
rect 197636 265202 197688 265208
rect 196532 265192 196584 265198
rect 196532 265134 196584 265140
rect 196440 147620 196492 147626
rect 196440 147562 196492 147568
rect 196544 147558 196572 265134
rect 196716 261180 196768 261186
rect 196716 261122 196768 261128
rect 196624 259684 196676 259690
rect 196624 259626 196676 259632
rect 196532 147552 196584 147558
rect 196532 147494 196584 147500
rect 196636 143410 196664 259626
rect 196728 146946 196756 261122
rect 197544 199096 197596 199102
rect 197544 199038 197596 199044
rect 197360 197124 197412 197130
rect 197360 197066 197412 197072
rect 196808 192432 196860 192438
rect 196808 192374 196860 192380
rect 196716 146940 196768 146946
rect 196716 146882 196768 146888
rect 196624 143404 196676 143410
rect 196624 143346 196676 143352
rect 196348 141840 196400 141846
rect 196348 141782 196400 141788
rect 196624 140480 196676 140486
rect 196624 140422 196676 140428
rect 196440 140072 196492 140078
rect 196440 140014 196492 140020
rect 196256 78668 196308 78674
rect 196256 78610 196308 78616
rect 196268 78130 196296 78610
rect 196256 78124 196308 78130
rect 196256 78066 196308 78072
rect 196452 71602 196480 140014
rect 196530 138000 196586 138009
rect 196530 137935 196586 137944
rect 196440 71596 196492 71602
rect 196440 71538 196492 71544
rect 196544 70242 196572 137935
rect 196636 78674 196664 140422
rect 196820 79218 196848 192374
rect 196992 147212 197044 147218
rect 196992 147154 197044 147160
rect 196900 144900 196952 144906
rect 196900 144842 196952 144848
rect 196808 79212 196860 79218
rect 196808 79154 196860 79160
rect 196624 78668 196676 78674
rect 196624 78610 196676 78616
rect 196912 71466 196940 144842
rect 197004 74322 197032 147154
rect 197084 147076 197136 147082
rect 197084 147018 197136 147024
rect 197096 81025 197124 147018
rect 197082 81016 197138 81025
rect 197082 80951 197138 80960
rect 196992 74316 197044 74322
rect 196992 74258 197044 74264
rect 196900 71460 196952 71466
rect 196900 71402 196952 71408
rect 196624 71120 196676 71126
rect 196624 71062 196676 71068
rect 196532 70236 196584 70242
rect 196532 70178 196584 70184
rect 196162 66736 196218 66745
rect 196162 66671 196218 66680
rect 196084 64846 196204 64874
rect 196070 62112 196126 62121
rect 196070 62047 196126 62056
rect 196084 61946 196112 62047
rect 196072 61940 196124 61946
rect 196072 61882 196124 61888
rect 196084 60790 196112 61882
rect 196072 60784 196124 60790
rect 196072 60726 196124 60732
rect 196176 58721 196204 64846
rect 196162 58712 196218 58721
rect 196162 58647 196218 58656
rect 195978 49464 196034 49473
rect 195978 49399 196034 49408
rect 195992 49065 196020 49399
rect 195978 49056 196034 49065
rect 195978 48991 196034 49000
rect 194598 47696 194654 47705
rect 194598 47631 194654 47640
rect 194598 44976 194654 44985
rect 194598 44911 194654 44920
rect 194612 16574 194640 44911
rect 194612 16546 195192 16574
rect 193864 3596 193916 3602
rect 193864 3538 193916 3544
rect 193784 3454 194456 3482
rect 194428 480 194456 3454
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196636 4146 196664 71062
rect 197372 62234 197400 197066
rect 197452 196920 197504 196926
rect 197452 196862 197504 196868
rect 197280 62206 197400 62234
rect 197280 61282 197308 62206
rect 197360 62076 197412 62082
rect 197360 62018 197412 62024
rect 197372 61470 197400 62018
rect 197360 61464 197412 61470
rect 197360 61406 197412 61412
rect 197280 61254 197400 61282
rect 197372 56273 197400 61254
rect 197358 56264 197414 56273
rect 197358 56199 197414 56208
rect 197360 55956 197412 55962
rect 197360 55898 197412 55904
rect 197372 16574 197400 55898
rect 197464 55185 197492 196862
rect 197556 62082 197584 199038
rect 197648 143002 197676 265202
rect 197912 265056 197964 265062
rect 197912 264998 197964 265004
rect 197820 261384 197872 261390
rect 197820 261326 197872 261332
rect 197728 259548 197780 259554
rect 197728 259490 197780 259496
rect 197636 142996 197688 143002
rect 197636 142938 197688 142944
rect 197740 141778 197768 259490
rect 197832 143274 197860 261326
rect 197924 147490 197952 264998
rect 218072 263430 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 234632 278089 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700670 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 234618 278080 234674 278089
rect 234618 278015 234674 278024
rect 282932 263498 282960 702406
rect 299492 276729 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 700466 332548 703520
rect 348804 702434 348832 703520
rect 364996 702434 365024 703520
rect 347792 702406 348832 702434
rect 364352 702406 365024 702434
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 299478 276720 299534 276729
rect 299478 276655 299534 276664
rect 282920 263492 282972 263498
rect 282920 263434 282972 263440
rect 218060 263424 218112 263430
rect 218060 263366 218112 263372
rect 347792 262886 347820 702406
rect 364352 273970 364380 702406
rect 397472 699718 397500 703520
rect 413664 700398 413692 703520
rect 413652 700392 413704 700398
rect 413652 700334 413704 700340
rect 429856 699718 429884 703520
rect 396724 699712 396776 699718
rect 396724 699654 396776 699660
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 428464 699712 428516 699718
rect 428464 699654 428516 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 396736 284986 396764 699654
rect 396724 284980 396776 284986
rect 396724 284922 396776 284928
rect 428476 275330 428504 699654
rect 462332 287706 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 462320 287700 462372 287706
rect 462320 287642 462372 287648
rect 428464 275324 428516 275330
rect 428464 275266 428516 275272
rect 364340 273964 364392 273970
rect 364340 273906 364392 273912
rect 347780 262880 347832 262886
rect 477512 262857 477540 702406
rect 489184 700392 489236 700398
rect 489184 700334 489236 700340
rect 489196 283626 489224 700334
rect 489184 283620 489236 283626
rect 489184 283562 489236 283568
rect 494072 271182 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 527824 700392 527876 700398
rect 527824 700334 527876 700340
rect 498844 670744 498896 670750
rect 498844 670686 498896 670692
rect 494060 271176 494112 271182
rect 494060 271118 494112 271124
rect 498856 268394 498884 670686
rect 527836 269822 527864 700334
rect 543476 700330 543504 703520
rect 559668 700398 559696 703520
rect 559656 700392 559708 700398
rect 559656 700334 559708 700340
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 527824 269816 527876 269822
rect 527824 269758 527876 269764
rect 498844 268388 498896 268394
rect 498844 268330 498896 268336
rect 580276 263566 580304 365055
rect 580264 263560 580316 263566
rect 580264 263502 580316 263508
rect 580356 263084 580408 263090
rect 580356 263026 580408 263032
rect 347780 262822 347832 262828
rect 477498 262848 477554 262857
rect 477498 262783 477554 262792
rect 200580 261520 200632 261526
rect 200580 261462 200632 261468
rect 199292 261248 199344 261254
rect 199292 261190 199344 261196
rect 199200 260908 199252 260914
rect 199200 260850 199252 260856
rect 198096 198076 198148 198082
rect 198096 198018 198148 198024
rect 197912 147484 197964 147490
rect 197912 147426 197964 147432
rect 198108 146305 198136 198018
rect 199108 198008 199160 198014
rect 199108 197950 199160 197956
rect 198832 197056 198884 197062
rect 198832 196998 198884 197004
rect 198738 196888 198794 196897
rect 198738 196823 198794 196832
rect 198188 152924 198240 152930
rect 198188 152866 198240 152872
rect 198094 146296 198150 146305
rect 198094 146231 198150 146240
rect 198004 145852 198056 145858
rect 198004 145794 198056 145800
rect 197820 143268 197872 143274
rect 197820 143210 197872 143216
rect 197728 141772 197780 141778
rect 197728 141714 197780 141720
rect 198016 78985 198044 145794
rect 198094 137864 198150 137873
rect 198094 137799 198150 137808
rect 198002 78976 198058 78985
rect 198002 78911 198058 78920
rect 198108 73098 198136 137799
rect 198096 73092 198148 73098
rect 198096 73034 198148 73040
rect 198200 69970 198228 152866
rect 198464 148640 198516 148646
rect 198464 148582 198516 148588
rect 198280 147008 198332 147014
rect 198280 146950 198332 146956
rect 198292 74390 198320 146950
rect 198372 143336 198424 143342
rect 198372 143278 198424 143284
rect 198280 74384 198332 74390
rect 198280 74326 198332 74332
rect 198188 69964 198240 69970
rect 198188 69906 198240 69912
rect 197544 62076 197596 62082
rect 197544 62018 197596 62024
rect 197636 62008 197688 62014
rect 197636 61950 197688 61956
rect 197648 61402 197676 61950
rect 198384 61402 198412 143278
rect 198476 75886 198504 148582
rect 198464 75880 198516 75886
rect 198464 75822 198516 75828
rect 197636 61396 197688 61402
rect 197636 61338 197688 61344
rect 198372 61396 198424 61402
rect 198372 61338 198424 61344
rect 197450 55176 197506 55185
rect 197450 55111 197506 55120
rect 197464 54505 197492 55111
rect 197450 54496 197506 54505
rect 197450 54431 197506 54440
rect 198752 50969 198780 196823
rect 198844 57361 198872 196998
rect 199016 196784 199068 196790
rect 199016 196726 199068 196732
rect 198924 196716 198976 196722
rect 198924 196658 198976 196664
rect 198936 60625 198964 196658
rect 199028 61849 199056 196726
rect 199120 80889 199148 197950
rect 199212 146198 199240 260850
rect 199304 148374 199332 261190
rect 200488 261044 200540 261050
rect 200488 260986 200540 260992
rect 200302 200288 200358 200297
rect 200302 200223 200358 200232
rect 200118 196752 200174 196761
rect 200118 196687 200174 196696
rect 199568 152856 199620 152862
rect 199568 152798 199620 152804
rect 199476 148504 199528 148510
rect 199476 148446 199528 148452
rect 199384 148436 199436 148442
rect 199384 148378 199436 148384
rect 199292 148368 199344 148374
rect 199292 148310 199344 148316
rect 199200 146192 199252 146198
rect 199200 146134 199252 146140
rect 199106 80880 199162 80889
rect 199106 80815 199162 80824
rect 199396 70038 199424 148378
rect 199488 72962 199516 148446
rect 199476 72956 199528 72962
rect 199476 72898 199528 72904
rect 199580 70174 199608 152798
rect 199660 148776 199712 148782
rect 199660 148718 199712 148724
rect 199568 70168 199620 70174
rect 199568 70110 199620 70116
rect 199672 70106 199700 148718
rect 199660 70100 199712 70106
rect 199660 70042 199712 70048
rect 199384 70032 199436 70038
rect 199384 69974 199436 69980
rect 199382 68912 199438 68921
rect 199382 68847 199384 68856
rect 199436 68847 199438 68856
rect 199384 68818 199436 68824
rect 199396 67658 199424 68818
rect 199384 67652 199436 67658
rect 199384 67594 199436 67600
rect 199014 61840 199070 61849
rect 199014 61775 199070 61784
rect 199028 61441 199056 61775
rect 199014 61432 199070 61441
rect 199014 61367 199070 61376
rect 198922 60616 198978 60625
rect 198922 60551 198978 60560
rect 198830 57352 198886 57361
rect 198830 57287 198886 57296
rect 198738 50960 198794 50969
rect 198738 50895 198794 50904
rect 199566 50960 199622 50969
rect 199566 50895 199622 50904
rect 199580 50289 199608 50895
rect 199566 50280 199622 50289
rect 199566 50215 199622 50224
rect 200132 49609 200160 196687
rect 200210 196616 200266 196625
rect 200210 196551 200266 196560
rect 200224 53825 200252 196551
rect 200316 63481 200344 200223
rect 200396 199368 200448 199374
rect 200396 199310 200448 199316
rect 200408 67590 200436 199310
rect 200500 145586 200528 260986
rect 200592 147354 200620 261462
rect 471244 261452 471296 261458
rect 471244 261394 471296 261400
rect 203248 259820 203300 259826
rect 203248 259762 203300 259768
rect 201774 200152 201830 200161
rect 201774 200087 201830 200096
rect 201684 199300 201736 199306
rect 201684 199242 201736 199248
rect 201040 198756 201092 198762
rect 201040 198698 201092 198704
rect 200672 152788 200724 152794
rect 200672 152730 200724 152736
rect 200580 147348 200632 147354
rect 200580 147290 200632 147296
rect 200488 145580 200540 145586
rect 200488 145522 200540 145528
rect 200396 67584 200448 67590
rect 200396 67526 200448 67532
rect 200302 63472 200358 63481
rect 200302 63407 200358 63416
rect 200210 53816 200266 53825
rect 200210 53751 200266 53760
rect 200118 49600 200174 49609
rect 200118 49535 200174 49544
rect 200684 44169 200712 152730
rect 200948 148912 201000 148918
rect 200948 148854 201000 148860
rect 200856 148844 200908 148850
rect 200856 148786 200908 148792
rect 200764 148572 200816 148578
rect 200764 148514 200816 148520
rect 200776 80986 200804 148514
rect 200764 80980 200816 80986
rect 200764 80922 200816 80928
rect 200868 69902 200896 148786
rect 200960 74526 200988 148854
rect 201052 147801 201080 198698
rect 201592 192364 201644 192370
rect 201592 192306 201644 192312
rect 201038 147792 201094 147801
rect 201038 147727 201094 147736
rect 201500 75540 201552 75546
rect 201500 75482 201552 75488
rect 200948 74520 201000 74526
rect 200948 74462 201000 74468
rect 200856 69896 200908 69902
rect 200856 69838 200908 69844
rect 200762 69592 200818 69601
rect 200762 69527 200818 69536
rect 200670 44160 200726 44169
rect 200670 44095 200726 44104
rect 198740 31408 198792 31414
rect 198740 31350 198792 31356
rect 197372 16546 197952 16574
rect 196624 4140 196676 4146
rect 196624 4082 196676 4088
rect 196808 3596 196860 3602
rect 196808 3538 196860 3544
rect 196820 480 196848 3538
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 31350
rect 200304 4140 200356 4146
rect 200304 4082 200356 4088
rect 200316 480 200344 4082
rect 200776 3194 200804 69527
rect 201408 67584 201460 67590
rect 201408 67526 201460 67532
rect 201420 66910 201448 67526
rect 201408 66904 201460 66910
rect 201408 66846 201460 66852
rect 201406 63472 201462 63481
rect 201406 63407 201462 63416
rect 201420 62937 201448 63407
rect 201406 62928 201462 62937
rect 201406 62863 201462 62872
rect 201406 53816 201462 53825
rect 201406 53751 201462 53760
rect 201420 53145 201448 53751
rect 201406 53136 201462 53145
rect 201406 53071 201462 53080
rect 201406 49600 201462 49609
rect 201406 49535 201462 49544
rect 201420 48929 201448 49535
rect 201406 48920 201462 48929
rect 201406 48855 201462 48864
rect 201512 11694 201540 75482
rect 201604 60058 201632 192306
rect 201696 64874 201724 199242
rect 201788 69834 201816 200087
rect 203156 193928 203208 193934
rect 203156 193870 203208 193876
rect 201868 193860 201920 193866
rect 201868 193802 201920 193808
rect 201880 79014 201908 193802
rect 202880 192840 202932 192846
rect 202880 192782 202932 192788
rect 202420 192704 202472 192710
rect 202420 192646 202472 192652
rect 202328 155236 202380 155242
rect 202328 155178 202380 155184
rect 202052 152652 202104 152658
rect 202052 152594 202104 152600
rect 201960 148708 202012 148714
rect 201960 148650 202012 148656
rect 201868 79008 201920 79014
rect 201868 78950 201920 78956
rect 201776 69828 201828 69834
rect 201776 69770 201828 69776
rect 201696 64846 201908 64874
rect 201604 60030 201816 60058
rect 201684 55208 201736 55214
rect 201682 55176 201684 55185
rect 201736 55176 201738 55185
rect 201682 55111 201738 55120
rect 201788 52465 201816 60030
rect 201880 59265 201908 64846
rect 201866 59256 201922 59265
rect 201866 59191 201922 59200
rect 201972 56545 202000 148650
rect 202064 69018 202092 152594
rect 202236 152584 202288 152590
rect 202236 152526 202288 152532
rect 202144 152516 202196 152522
rect 202144 152458 202196 152464
rect 202156 70378 202184 152458
rect 202144 70372 202196 70378
rect 202144 70314 202196 70320
rect 202248 70310 202276 152526
rect 202340 73166 202368 155178
rect 202328 73160 202380 73166
rect 202328 73102 202380 73108
rect 202432 72894 202460 192646
rect 202420 72888 202472 72894
rect 202420 72830 202472 72836
rect 202432 72486 202460 72830
rect 202420 72480 202472 72486
rect 202420 72422 202472 72428
rect 202236 70304 202288 70310
rect 202236 70246 202288 70252
rect 202788 69828 202840 69834
rect 202788 69770 202840 69776
rect 202800 69698 202828 69770
rect 202788 69692 202840 69698
rect 202788 69634 202840 69640
rect 202052 69012 202104 69018
rect 202052 68954 202104 68960
rect 202786 59256 202842 59265
rect 202786 59191 202842 59200
rect 202800 58585 202828 59191
rect 202786 58576 202842 58585
rect 202786 58511 202842 58520
rect 201958 56536 202014 56545
rect 201958 56471 202014 56480
rect 202786 56536 202842 56545
rect 202786 56471 202842 56480
rect 202800 56137 202828 56471
rect 202786 56128 202842 56137
rect 202786 56063 202842 56072
rect 202788 55208 202840 55214
rect 202788 55150 202840 55156
rect 202800 53854 202828 55150
rect 202788 53848 202840 53854
rect 202788 53790 202840 53796
rect 201774 52456 201830 52465
rect 201774 52391 201830 52400
rect 202786 52456 202842 52465
rect 202786 52391 202842 52400
rect 202800 51785 202828 52391
rect 202786 51776 202842 51785
rect 202786 51711 202842 51720
rect 201592 47796 201644 47802
rect 201592 47738 201644 47744
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 47738
rect 202892 44033 202920 192782
rect 203064 192772 203116 192778
rect 203064 192714 203116 192720
rect 202972 192636 203024 192642
rect 202972 192578 203024 192584
rect 202984 52426 203012 192578
rect 203076 64870 203104 192714
rect 203168 77353 203196 193870
rect 203260 149870 203288 259762
rect 471256 206990 471284 261394
rect 472624 259480 472676 259486
rect 472624 259422 472676 259428
rect 472636 245614 472664 259422
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 472624 245608 472676 245614
rect 580172 245608 580224 245614
rect 472624 245550 472676 245556
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580368 219065 580396 263026
rect 580448 262948 580500 262954
rect 580448 262890 580500 262896
rect 580460 232393 580488 262890
rect 580446 232384 580502 232393
rect 580446 232319 580502 232328
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 471244 206984 471296 206990
rect 471244 206926 471296 206932
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 205730 193080 205786 193089
rect 205730 193015 205786 193024
rect 204258 192672 204314 192681
rect 204258 192607 204314 192616
rect 203340 155440 203392 155446
rect 203340 155382 203392 155388
rect 203248 149864 203300 149870
rect 203248 149806 203300 149812
rect 203154 77344 203210 77353
rect 203154 77279 203210 77288
rect 203064 64864 203116 64870
rect 203064 64806 203116 64812
rect 203076 64190 203104 64806
rect 203064 64184 203116 64190
rect 203064 64126 203116 64132
rect 202972 52420 203024 52426
rect 202972 52362 203024 52368
rect 203064 51060 203116 51066
rect 203064 51002 203116 51008
rect 203076 50969 203104 51002
rect 203062 50960 203118 50969
rect 203062 50895 203118 50904
rect 203352 48249 203380 155382
rect 203524 155372 203576 155378
rect 203524 155314 203576 155320
rect 203432 155304 203484 155310
rect 203432 155246 203484 155252
rect 203444 57934 203472 155246
rect 203536 71534 203564 155314
rect 203800 152720 203852 152726
rect 203800 152662 203852 152668
rect 203708 150136 203760 150142
rect 203708 150078 203760 150084
rect 203616 150000 203668 150006
rect 203616 149942 203668 149948
rect 203524 71528 203576 71534
rect 203524 71470 203576 71476
rect 203628 68241 203656 149942
rect 203720 78305 203748 150078
rect 203706 78296 203762 78305
rect 203706 78231 203762 78240
rect 203708 76560 203760 76566
rect 203708 76502 203760 76508
rect 203614 68232 203670 68241
rect 203614 68167 203670 68176
rect 203432 57928 203484 57934
rect 203432 57870 203484 57876
rect 203338 48240 203394 48249
rect 203338 48175 203394 48184
rect 202878 44024 202934 44033
rect 202878 43959 202934 43968
rect 202892 43489 202920 43959
rect 202878 43480 202934 43489
rect 202878 43415 202934 43424
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 200764 3188 200816 3194
rect 200764 3130 200816 3136
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 203720 3670 203748 76502
rect 203812 53786 203840 152662
rect 204166 78024 204222 78033
rect 204166 77959 204222 77968
rect 204180 77353 204208 77959
rect 204166 77344 204222 77353
rect 204166 77279 204222 77288
rect 204168 57928 204220 57934
rect 204168 57870 204220 57876
rect 204180 57254 204208 57870
rect 204168 57248 204220 57254
rect 204168 57190 204220 57196
rect 204272 56001 204300 192607
rect 205640 192568 205692 192574
rect 205640 192510 205692 192516
rect 204352 150068 204404 150074
rect 204352 150010 204404 150016
rect 204258 55992 204314 56001
rect 204258 55927 204314 55936
rect 204260 55888 204312 55894
rect 204260 55830 204312 55836
rect 203800 53780 203852 53786
rect 203800 53722 203852 53728
rect 203812 53106 203840 53722
rect 203800 53100 203852 53106
rect 203800 53042 203852 53048
rect 204168 52420 204220 52426
rect 204168 52362 204220 52368
rect 204180 51746 204208 52362
rect 204168 51740 204220 51746
rect 204168 51682 204220 51688
rect 204168 51060 204220 51066
rect 204168 51002 204220 51008
rect 204180 49774 204208 51002
rect 204168 49768 204220 49774
rect 204168 49710 204220 49716
rect 204166 48240 204222 48249
rect 204166 48175 204222 48184
rect 204180 47569 204208 48175
rect 204166 47560 204222 47569
rect 204166 47495 204222 47504
rect 204272 16574 204300 55830
rect 204364 46918 204392 150010
rect 204536 149932 204588 149938
rect 204536 149874 204588 149880
rect 204444 149728 204496 149734
rect 204444 149670 204496 149676
rect 204456 71738 204484 149670
rect 204548 72350 204576 149874
rect 204628 149796 204680 149802
rect 204628 149738 204680 149744
rect 204640 76673 204668 149738
rect 204626 76664 204682 76673
rect 204626 76599 204682 76608
rect 205652 73137 205680 192510
rect 205744 75070 205772 193015
rect 205914 192944 205970 192953
rect 205914 192879 205970 192888
rect 206100 192908 206152 192914
rect 205822 192536 205878 192545
rect 205822 192471 205878 192480
rect 205836 78402 205864 192471
rect 205824 78396 205876 78402
rect 205824 78338 205876 78344
rect 205824 77240 205876 77246
rect 205824 77182 205876 77188
rect 205836 76566 205864 77182
rect 205928 77042 205956 192879
rect 206100 192850 206152 192856
rect 206006 192808 206062 192817
rect 206006 192743 206062 192752
rect 205916 77036 205968 77042
rect 205916 76978 205968 76984
rect 205914 76936 205970 76945
rect 206020 76922 206048 192743
rect 206112 77246 206140 192850
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 206192 192500 206244 192506
rect 580170 192471 580226 192480
rect 206192 192442 206244 192448
rect 206204 80918 206232 192442
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580354 152688 580410 152697
rect 580354 152623 580410 152632
rect 580264 146328 580316 146334
rect 580264 146270 580316 146276
rect 327724 140888 327776 140894
rect 327724 140830 327776 140836
rect 289082 139632 289138 139641
rect 289082 139567 289138 139576
rect 206192 80912 206244 80918
rect 206192 80854 206244 80860
rect 234620 80912 234672 80918
rect 234620 80854 234672 80860
rect 206192 78396 206244 78402
rect 206192 78338 206244 78344
rect 206100 77240 206152 77246
rect 206100 77182 206152 77188
rect 205970 76894 206048 76922
rect 205914 76871 205970 76880
rect 205824 76560 205876 76566
rect 205928 76537 205956 76871
rect 205824 76502 205876 76508
rect 205914 76528 205970 76537
rect 205914 76463 205970 76472
rect 206204 75721 206232 78338
rect 211802 76800 211858 76809
rect 211802 76735 211858 76744
rect 206190 75712 206246 75721
rect 206190 75647 206246 75656
rect 206558 75712 206614 75721
rect 206558 75647 206614 75656
rect 206572 75177 206600 75647
rect 206558 75168 206614 75177
rect 206558 75103 206614 75112
rect 205732 75064 205784 75070
rect 205732 75006 205784 75012
rect 205638 73128 205694 73137
rect 205638 73063 205694 73072
rect 206284 73092 206336 73098
rect 205652 72457 205680 73063
rect 206284 73034 206336 73040
rect 205638 72448 205694 72457
rect 205638 72383 205694 72392
rect 204536 72344 204588 72350
rect 204536 72286 204588 72292
rect 204444 71732 204496 71738
rect 204444 71674 204496 71680
rect 204456 71126 204484 71674
rect 204444 71120 204496 71126
rect 204444 71062 204496 71068
rect 204352 46912 204404 46918
rect 204352 46854 204404 46860
rect 204720 46912 204772 46918
rect 204720 46854 204772 46860
rect 204732 46238 204760 46854
rect 204720 46232 204772 46238
rect 204720 46174 204772 46180
rect 205640 40996 205692 41002
rect 205640 40938 205692 40944
rect 205652 16574 205680 40938
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 203708 3664 203760 3670
rect 203708 3606 203760 3612
rect 203892 3188 203944 3194
rect 203892 3130 203944 3136
rect 203904 480 203932 3130
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 206296 3602 206324 73034
rect 207020 65612 207072 65618
rect 207020 65554 207072 65560
rect 206284 3596 206336 3602
rect 206284 3538 206336 3544
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207032 354 207060 65554
rect 209872 54596 209924 54602
rect 209872 54538 209924 54544
rect 208400 47728 208452 47734
rect 208400 47670 208452 47676
rect 208412 16574 208440 47670
rect 208412 16546 208624 16574
rect 208596 480 208624 16546
rect 209884 6914 209912 54538
rect 209792 6886 209912 6914
rect 209792 480 209820 6886
rect 211816 3806 211844 76735
rect 216680 75472 216732 75478
rect 216680 75414 216732 75420
rect 213918 67144 213974 67153
rect 213918 67079 213974 67088
rect 212538 32464 212594 32473
rect 212538 32399 212594 32408
rect 212552 16574 212580 32399
rect 213932 16574 213960 67079
rect 215300 53236 215352 53242
rect 215300 53178 215352 53184
rect 212552 16546 213408 16574
rect 213932 16546 214512 16574
rect 210976 3800 211028 3806
rect 210976 3742 211028 3748
rect 211804 3800 211856 3806
rect 211804 3742 211856 3748
rect 210988 480 211016 3742
rect 212172 3732 212224 3738
rect 212172 3674 212224 3680
rect 212184 480 212212 3674
rect 213380 480 213408 16546
rect 214484 480 214512 16546
rect 207358 354 207470 480
rect 207032 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 53178
rect 216692 16574 216720 75414
rect 218060 71120 218112 71126
rect 218060 71062 218112 71068
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 480 218100 71062
rect 220820 68468 220872 68474
rect 220820 68410 220872 68416
rect 218152 50516 218204 50522
rect 218152 50458 218204 50464
rect 218164 16574 218192 50458
rect 219440 23044 219492 23050
rect 219440 22986 219492 22992
rect 219452 16574 219480 22986
rect 220832 16574 220860 68410
rect 224960 64320 225012 64326
rect 224960 64262 225012 64268
rect 223580 60240 223632 60246
rect 223580 60182 223632 60188
rect 222200 49156 222252 49162
rect 222200 49098 222252 49104
rect 222212 16574 222240 49098
rect 218164 16546 219296 16574
rect 219452 16546 220032 16574
rect 220832 16546 221136 16574
rect 222212 16546 222792 16574
rect 219268 480 219296 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 16546
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 16546
rect 222764 480 222792 16546
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 60182
rect 224972 16574 225000 64262
rect 227718 63336 227774 63345
rect 227718 63271 227774 63280
rect 226340 36780 226392 36786
rect 226340 36722 226392 36728
rect 224972 16546 225184 16574
rect 225156 480 225184 16546
rect 226352 480 226380 36722
rect 227732 16574 227760 63271
rect 231858 61704 231914 61713
rect 231858 61639 231914 61648
rect 230478 42120 230534 42129
rect 230478 42055 230534 42064
rect 229098 18592 229154 18601
rect 229098 18527 229154 18536
rect 229112 16574 229140 18527
rect 230492 16574 230520 42055
rect 227732 16546 228312 16574
rect 229112 16546 229416 16574
rect 230492 16546 231072 16574
rect 227536 7812 227588 7818
rect 227536 7754 227588 7760
rect 227548 480 227576 7754
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 229388 354 229416 16546
rect 231044 480 231072 16546
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 228702 -960 228814 326
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 231872 354 231900 61639
rect 233240 57316 233292 57322
rect 233240 57258 233292 57264
rect 233252 16574 233280 57258
rect 233252 16546 233464 16574
rect 233436 480 233464 16546
rect 234632 3806 234660 80854
rect 252560 80844 252612 80850
rect 252560 80786 252612 80792
rect 238760 80096 238812 80102
rect 238760 80038 238812 80044
rect 237380 74248 237432 74254
rect 237380 74190 237432 74196
rect 236000 46436 236052 46442
rect 236000 46378 236052 46384
rect 236012 16574 236040 46378
rect 237392 16574 237420 74190
rect 238772 16574 238800 80038
rect 247682 76664 247738 76673
rect 247682 76599 247738 76608
rect 242898 67280 242954 67289
rect 242898 67215 242954 67224
rect 241520 17536 241572 17542
rect 241520 17478 241572 17484
rect 241532 16574 241560 17478
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 241532 16546 241744 16574
rect 234712 9308 234764 9314
rect 234712 9250 234764 9256
rect 234620 3800 234672 3806
rect 234620 3742 234672 3748
rect 234724 3482 234752 9250
rect 235816 3800 235868 3806
rect 235816 3742 235868 3748
rect 234632 3454 234752 3482
rect 234632 480 234660 3454
rect 235828 480 235856 3742
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 240508 3664 240560 3670
rect 240508 3606 240560 3612
rect 240520 480 240548 3606
rect 241716 480 241744 16546
rect 242912 480 242940 67215
rect 245660 60172 245712 60178
rect 245660 60114 245712 60120
rect 242992 28552 243044 28558
rect 242992 28494 243044 28500
rect 243004 16574 243032 28494
rect 245672 16574 245700 60114
rect 243004 16546 244136 16574
rect 245672 16546 245976 16574
rect 244108 480 244136 16546
rect 245200 11960 245252 11966
rect 245200 11902 245252 11908
rect 245212 480 245240 11902
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247592 3732 247644 3738
rect 247592 3674 247644 3680
rect 247604 480 247632 3674
rect 247696 3670 247724 76599
rect 248420 73840 248472 73846
rect 248420 73782 248472 73788
rect 247684 3664 247736 3670
rect 247684 3606 247736 3612
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 73782
rect 249798 44840 249854 44849
rect 249798 44775 249854 44784
rect 249812 16574 249840 44775
rect 251180 39636 251232 39642
rect 251180 39578 251232 39584
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 480 251220 39578
rect 251272 34060 251324 34066
rect 251272 34002 251324 34008
rect 251284 16574 251312 34002
rect 252572 16574 252600 80786
rect 270500 80776 270552 80782
rect 270500 80718 270552 80724
rect 253204 78328 253256 78334
rect 253204 78270 253256 78276
rect 253216 73846 253244 78270
rect 269762 78024 269818 78033
rect 269762 77959 269818 77968
rect 260840 76764 260892 76770
rect 260840 76706 260892 76712
rect 255320 74180 255372 74186
rect 255320 74122 255372 74128
rect 253204 73840 253256 73846
rect 253204 73782 253256 73788
rect 255332 16574 255360 74122
rect 256700 64252 256752 64258
rect 256700 64194 256752 64200
rect 251284 16546 252416 16574
rect 252572 16546 253520 16574
rect 255332 16546 255912 16574
rect 252388 480 252416 16546
rect 253492 480 253520 16546
rect 254676 3664 254728 3670
rect 254676 3606 254728 3612
rect 254688 480 254716 3606
rect 255884 480 255912 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 354 256740 64194
rect 259460 50448 259512 50454
rect 259460 50390 259512 50396
rect 259472 11694 259500 50390
rect 260852 16574 260880 76706
rect 269120 74452 269172 74458
rect 269120 74394 269172 74400
rect 261484 73908 261536 73914
rect 261484 73850 261536 73856
rect 260852 16546 261432 16574
rect 259552 16176 259604 16182
rect 259552 16118 259604 16124
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 258264 10600 258316 10606
rect 258264 10542 258316 10548
rect 258276 480 258304 10542
rect 259564 6914 259592 16118
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261404 3482 261432 16546
rect 261496 3670 261524 73850
rect 263598 57760 263654 57769
rect 263598 57695 263654 57704
rect 263612 16574 263640 57695
rect 267738 40624 267794 40633
rect 267738 40559 267794 40568
rect 264978 26888 265034 26897
rect 264978 26823 265034 26832
rect 263612 16546 264192 16574
rect 261484 3664 261536 3670
rect 261484 3606 261536 3612
rect 262956 3664 263008 3670
rect 262956 3606 263008 3612
rect 261404 3454 261800 3482
rect 261772 480 261800 3454
rect 262968 480 262996 3606
rect 264164 480 264192 16546
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 26823
rect 266544 5024 266596 5030
rect 266544 4966 266596 4972
rect 266556 480 266584 4966
rect 267752 480 267780 40559
rect 267832 32632 267884 32638
rect 267832 32574 267884 32580
rect 267844 16574 267872 32574
rect 269132 16574 269160 74394
rect 269776 73914 269804 77959
rect 269764 73908 269816 73914
rect 269764 73850 269816 73856
rect 270512 16574 270540 80718
rect 288440 78940 288492 78946
rect 288440 78882 288492 78888
rect 287702 77888 287758 77897
rect 287702 77823 287758 77832
rect 284300 74112 284352 74118
rect 284300 74054 284352 74060
rect 274638 65920 274694 65929
rect 274638 65855 274694 65864
rect 273260 20256 273312 20262
rect 273260 20198 273312 20204
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 272432 14748 272484 14754
rect 272432 14690 272484 14696
rect 272444 480 272472 14690
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 20198
rect 274652 16574 274680 65855
rect 277398 63200 277454 63209
rect 277398 63135 277454 63144
rect 275284 46368 275336 46374
rect 275284 46310 275336 46316
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 275296 3398 275324 46310
rect 277412 16574 277440 63135
rect 281538 58984 281594 58993
rect 281538 58919 281594 58928
rect 278780 25832 278832 25838
rect 278780 25774 278832 25780
rect 278792 16574 278820 25774
rect 280160 20188 280212 20194
rect 280160 20130 280212 20136
rect 280172 16574 280200 20130
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 276020 13388 276072 13394
rect 276020 13330 276072 13336
rect 275284 3392 275336 3398
rect 275284 3334 275336 3340
rect 276032 480 276060 13330
rect 277124 3392 277176 3398
rect 277124 3334 277176 3340
rect 277136 480 277164 3334
rect 278332 480 278360 16546
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 58919
rect 282920 24336 282972 24342
rect 282920 24278 282972 24284
rect 282932 16574 282960 24278
rect 282932 16546 283144 16574
rect 283116 480 283144 16546
rect 284312 480 284340 74054
rect 284390 53408 284446 53417
rect 284390 53343 284446 53352
rect 284404 16574 284432 53343
rect 285680 49088 285732 49094
rect 285680 49030 285732 49036
rect 285692 16574 285720 49030
rect 287716 19990 287744 77823
rect 287060 19984 287112 19990
rect 287060 19926 287112 19932
rect 287704 19984 287756 19990
rect 287704 19926 287756 19932
rect 287072 16574 287100 19926
rect 288452 16574 288480 78882
rect 289096 20670 289124 139567
rect 306380 79416 306432 79422
rect 306380 79358 306432 79364
rect 289820 76016 289872 76022
rect 289820 75958 289872 75964
rect 289084 20664 289136 20670
rect 289084 20606 289136 20612
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 354 284984 16546
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 75958
rect 296720 75948 296772 75954
rect 296720 75890 296772 75896
rect 295338 67008 295394 67017
rect 295338 66943 295394 66952
rect 292578 63064 292634 63073
rect 292578 62999 292634 63008
rect 291200 20120 291252 20126
rect 291200 20062 291252 20068
rect 291212 16574 291240 20062
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 292592 480 292620 62999
rect 292672 42356 292724 42362
rect 292672 42298 292724 42304
rect 292684 16574 292712 42298
rect 293960 38208 294012 38214
rect 293960 38150 294012 38156
rect 293972 16574 294000 38150
rect 295352 16574 295380 66943
rect 296732 16574 296760 75890
rect 297364 74044 297416 74050
rect 297364 73986 297416 73992
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 295352 16546 295656 16574
rect 296732 16546 297312 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297284 480 297312 16546
rect 297376 3194 297404 73986
rect 304998 73808 305054 73817
rect 304998 73743 305054 73752
rect 301502 72448 301558 72457
rect 301502 72383 301558 72392
rect 299480 60104 299532 60110
rect 299480 60046 299532 60052
rect 299492 3482 299520 60046
rect 299572 36712 299624 36718
rect 299572 36654 299624 36660
rect 299584 3670 299612 36654
rect 300860 18828 300912 18834
rect 300860 18770 300912 18776
rect 300872 6914 300900 18770
rect 301516 16574 301544 72383
rect 302240 68400 302292 68406
rect 302240 68342 302292 68348
rect 302252 16574 302280 68342
rect 303620 31340 303672 31346
rect 303620 31282 303672 31288
rect 303632 16574 303660 31282
rect 305012 16574 305040 73743
rect 301516 16546 301636 16574
rect 302252 16546 303200 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 300872 6886 301544 6914
rect 299572 3664 299624 3670
rect 299572 3606 299624 3612
rect 300768 3664 300820 3670
rect 300768 3606 300820 3612
rect 299492 3454 299704 3482
rect 297364 3188 297416 3194
rect 297364 3130 297416 3136
rect 298468 3188 298520 3194
rect 298468 3130 298520 3136
rect 298480 480 298508 3130
rect 299676 480 299704 3454
rect 300780 480 300808 3606
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 6886
rect 301608 4146 301636 16546
rect 301596 4140 301648 4146
rect 301596 4082 301648 4088
rect 303172 480 303200 16546
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306392 354 306420 79358
rect 324320 79348 324372 79354
rect 324320 79290 324372 79296
rect 311164 72820 311216 72826
rect 311164 72762 311216 72768
rect 309138 61568 309194 61577
rect 309138 61503 309194 61512
rect 309152 16574 309180 61503
rect 310520 35488 310572 35494
rect 310520 35430 310572 35436
rect 310532 16574 310560 35430
rect 309152 16546 309824 16574
rect 310532 16546 311112 16574
rect 307944 10532 307996 10538
rect 307944 10474 307996 10480
rect 307956 480 307984 10474
rect 309048 4140 309100 4146
rect 309048 4082 309100 4088
rect 309060 480 309088 4082
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311084 3482 311112 16546
rect 311176 3670 311204 72762
rect 318800 72752 318852 72758
rect 318800 72694 318852 72700
rect 313278 57624 313334 57633
rect 313278 57559 313334 57568
rect 313292 16574 313320 57559
rect 315304 43580 315356 43586
rect 315304 43522 315356 43528
rect 313292 16546 313872 16574
rect 311164 3664 311216 3670
rect 311164 3606 311216 3612
rect 312636 3664 312688 3670
rect 312636 3606 312688 3612
rect 311084 3454 311480 3482
rect 311452 480 311480 3454
rect 312648 480 312676 3606
rect 313844 480 313872 16546
rect 314660 14680 314712 14686
rect 314660 14622 314712 14628
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 14622
rect 315316 4146 315344 43522
rect 317420 40928 317472 40934
rect 317420 40870 317472 40876
rect 317432 16574 317460 40870
rect 318812 16574 318840 72694
rect 320180 51808 320232 51814
rect 320180 51750 320232 51756
rect 320192 16574 320220 51750
rect 321560 29912 321612 29918
rect 321560 29854 321612 29860
rect 321572 16574 321600 29854
rect 322940 21616 322992 21622
rect 322940 21558 322992 21564
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316224 6452 316276 6458
rect 316224 6394 316276 6400
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 316236 480 316264 6394
rect 317328 4140 317380 4146
rect 317328 4082 317380 4088
rect 317340 480 317368 4082
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 21558
rect 324332 3210 324360 79290
rect 327736 73166 327764 140830
rect 464344 140820 464396 140826
rect 464344 140762 464396 140768
rect 464356 86970 464384 140762
rect 576122 139496 576178 139505
rect 576122 139431 576178 139440
rect 464344 86964 464396 86970
rect 464344 86906 464396 86912
rect 523130 80880 523186 80889
rect 523130 80815 523186 80824
rect 358820 80708 358872 80714
rect 358820 80650 358872 80656
rect 337384 78260 337436 78266
rect 337384 78202 337436 78208
rect 327724 73160 327776 73166
rect 327724 73102 327776 73108
rect 324964 72684 325016 72690
rect 324964 72626 325016 72632
rect 324412 13320 324464 13326
rect 324412 13262 324464 13268
rect 324424 3398 324452 13262
rect 324976 4146 325004 72626
rect 332600 72616 332652 72622
rect 332600 72558 332652 72564
rect 327078 58848 327134 58857
rect 327078 58783 327134 58792
rect 327092 16574 327120 58783
rect 331218 54768 331274 54777
rect 331218 54703 331274 54712
rect 329840 21548 329892 21554
rect 329840 21490 329892 21496
rect 329852 16574 329880 21490
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 324964 4140 325016 4146
rect 324964 4082 325016 4088
rect 326804 4140 326856 4146
rect 326804 4082 326856 4088
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 326816 480 326844 4082
rect 328012 480 328040 16546
rect 329196 9240 329248 9246
rect 329196 9182 329248 9188
rect 329208 480 329236 9182
rect 330404 480 330432 16546
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 54703
rect 332612 3398 332640 72558
rect 332692 67720 332744 67726
rect 332692 67662 332744 67668
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 67662
rect 333980 53168 334032 53174
rect 333980 53110 334032 53116
rect 333992 16574 334020 53110
rect 337396 21486 337424 78202
rect 353300 76696 353352 76702
rect 353300 76638 353352 76644
rect 347780 73976 347832 73982
rect 347780 73918 347832 73924
rect 346400 65544 346452 65550
rect 346400 65486 346452 65492
rect 340880 62892 340932 62898
rect 340880 62834 340932 62840
rect 338118 50416 338174 50425
rect 338118 50351 338174 50360
rect 336740 21480 336792 21486
rect 336740 21422 336792 21428
rect 337384 21480 337436 21486
rect 337384 21422 337436 21428
rect 336752 16574 336780 21422
rect 338132 16574 338160 50351
rect 339500 28484 339552 28490
rect 339500 28426 339552 28432
rect 333992 16546 334664 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336278 11656 336334 11665
rect 336278 11591 336334 11600
rect 336292 480 336320 11591
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 28426
rect 340892 3398 340920 62834
rect 345020 60036 345072 60042
rect 345020 59978 345072 59984
rect 342260 35420 342312 35426
rect 342260 35362 342312 35368
rect 340972 31272 341024 31278
rect 340972 31214 341024 31220
rect 340880 3392 340932 3398
rect 340880 3334 340932 3340
rect 340984 480 341012 31214
rect 342272 16574 342300 35362
rect 343640 21412 343692 21418
rect 343640 21354 343692 21360
rect 343652 16574 343680 21354
rect 345032 16574 345060 59978
rect 346412 16574 346440 65486
rect 347792 16574 347820 73918
rect 349158 56400 349214 56409
rect 349158 56335 349214 56344
rect 349172 16574 349200 56335
rect 351920 38140 351972 38146
rect 351920 38082 351972 38088
rect 350540 22976 350592 22982
rect 350540 22918 350592 22924
rect 350552 16574 350580 22918
rect 351932 16574 351960 38082
rect 353312 16574 353340 76638
rect 354680 71052 354732 71058
rect 354680 70994 354732 71000
rect 354692 16574 354720 70994
rect 357440 62824 357492 62830
rect 357440 62766 357492 62772
rect 356058 49192 356114 49201
rect 356058 49127 356114 49136
rect 356072 16574 356100 49127
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 349172 16546 349292 16574
rect 350552 16546 351224 16574
rect 351932 16546 352880 16574
rect 353312 16546 353616 16574
rect 354692 16546 355272 16574
rect 356072 16546 356376 16574
rect 342168 3392 342220 3398
rect 342168 3334 342220 3340
rect 342180 480 342208 3334
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 344572 480 344600 16546
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349264 480 349292 16546
rect 350448 7744 350500 7750
rect 350448 7686 350500 7692
rect 350460 480 350488 7686
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352852 480 352880 16546
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355244 480 355272 16546
rect 356348 480 356376 16546
rect 357452 3398 357480 62766
rect 357532 32564 357584 32570
rect 357532 32506 357584 32512
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 32506
rect 358832 16574 358860 80650
rect 480260 78872 480312 78878
rect 382278 78840 382334 78849
rect 480260 78814 480312 78820
rect 382278 78775 382334 78784
rect 367100 76628 367152 76634
rect 367100 76570 367152 76576
rect 362958 65784 363014 65793
rect 362958 65719 363014 65728
rect 361580 39568 361632 39574
rect 361580 39510 361632 39516
rect 361592 16574 361620 39510
rect 362972 16574 363000 65719
rect 364982 57488 365038 57497
rect 364982 57423 365038 57432
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 16108 361172 16114
rect 361120 16050 361172 16056
rect 361132 480 361160 16050
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364616 16040 364668 16046
rect 364616 15982 364668 15988
rect 364628 480 364656 15982
rect 364996 3398 365024 57423
rect 367112 16574 367140 76570
rect 368480 72548 368532 72554
rect 368480 72490 368532 72496
rect 368492 16574 368520 72490
rect 376758 66872 376814 66881
rect 376758 66807 376814 66816
rect 369858 54632 369914 54641
rect 369858 54567 369914 54576
rect 369872 16574 369900 54567
rect 373998 47696 374054 47705
rect 373998 47631 374054 47640
rect 372620 20052 372672 20058
rect 372620 19994 372672 20000
rect 372632 16574 372660 19994
rect 367112 16546 367784 16574
rect 368492 16546 369440 16574
rect 369872 16546 370176 16574
rect 372632 16546 372936 16574
rect 365812 9172 365864 9178
rect 365812 9114 365864 9120
rect 364984 3392 365036 3398
rect 364984 3334 365036 3340
rect 365824 480 365852 9114
rect 367008 3392 367060 3398
rect 367008 3334 367060 3340
rect 367020 480 367048 3334
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371700 6384 371752 6390
rect 371700 6326 371752 6332
rect 371712 480 371740 6326
rect 372908 480 372936 16546
rect 374012 1170 374040 47631
rect 375380 29844 375432 29850
rect 375380 29786 375432 29792
rect 374092 27124 374144 27130
rect 374092 27066 374144 27072
rect 374104 3398 374132 27066
rect 375392 16574 375420 29786
rect 376772 16574 376800 66807
rect 380898 58712 380954 58721
rect 380898 58647 380954 58656
rect 379520 28416 379572 28422
rect 379520 28358 379572 28364
rect 375392 16546 376064 16574
rect 376772 16546 377720 16574
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 1142 374132 1170
rect 374104 480 374132 1142
rect 375300 480 375328 3334
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 378876 4956 378928 4962
rect 378876 4898 378928 4904
rect 378888 480 378916 4898
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379532 354 379560 28358
rect 380912 16574 380940 58647
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 3398 382320 78775
rect 436098 78704 436154 78713
rect 436098 78639 436154 78648
rect 400864 78192 400916 78198
rect 400864 78134 400916 78140
rect 389180 66972 389232 66978
rect 389180 66914 389232 66920
rect 382922 53272 382978 53281
rect 382922 53207 382978 53216
rect 382372 25764 382424 25770
rect 382372 25706 382424 25712
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 25706
rect 382936 4146 382964 53207
rect 387798 49056 387854 49065
rect 387798 48991 387854 49000
rect 386696 11892 386748 11898
rect 386696 11834 386748 11840
rect 385960 10464 386012 10470
rect 385960 10406 386012 10412
rect 382924 4140 382976 4146
rect 382924 4082 382976 4088
rect 384764 4140 384816 4146
rect 384764 4082 384816 4088
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 384776 480 384804 4082
rect 385972 480 386000 10406
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386708 354 386736 11834
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387812 354 387840 48991
rect 389192 16574 389220 66914
rect 394700 61464 394752 61470
rect 394700 61406 394752 61412
rect 390560 45008 390612 45014
rect 390560 44950 390612 44956
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3398 390600 44950
rect 391940 33992 391992 33998
rect 391940 33934 391992 33940
rect 391952 16574 391980 33934
rect 394712 16574 394740 61406
rect 396080 61396 396132 61402
rect 396080 61338 396132 61344
rect 391952 16546 392624 16574
rect 394712 16546 395384 16574
rect 390652 10396 390704 10402
rect 390652 10338 390704 10344
rect 390560 3392 390612 3398
rect 390560 3334 390612 3340
rect 390664 480 390692 10338
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394240 14612 394292 14618
rect 394240 14554 394292 14560
rect 394252 480 394280 14554
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 61338
rect 398838 56264 398894 56273
rect 398838 56199 398894 56208
rect 397736 15972 397788 15978
rect 397736 15914 397788 15920
rect 397748 480 397776 15914
rect 398852 3210 398880 56199
rect 398932 24268 398984 24274
rect 398932 24210 398984 24216
rect 398944 3398 398972 24210
rect 400876 15978 400904 78134
rect 429200 78124 429252 78130
rect 429200 78066 429252 78072
rect 415492 78056 415544 78062
rect 415492 77998 415544 78004
rect 412638 60072 412694 60081
rect 412638 60007 412694 60016
rect 401598 54496 401654 54505
rect 401598 54431 401654 54440
rect 401612 16574 401640 54431
rect 405738 51912 405794 51921
rect 405738 51847 405794 51856
rect 404360 43512 404412 43518
rect 404360 43454 404412 43460
rect 401612 16546 402560 16574
rect 400864 15972 400916 15978
rect 400864 15914 400916 15920
rect 400864 13252 400916 13258
rect 400864 13194 400916 13200
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 13194
rect 402532 480 402560 16546
rect 403624 3596 403676 3602
rect 403624 3538 403676 3544
rect 403636 480 403664 3538
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 43454
rect 405752 16574 405780 51847
rect 408500 43444 408552 43450
rect 408500 43386 408552 43392
rect 407120 27056 407172 27062
rect 407120 26998 407172 27004
rect 405752 16546 406056 16574
rect 406028 480 406056 16546
rect 407132 3602 407160 26998
rect 408512 16574 408540 43386
rect 410524 33924 410576 33930
rect 410524 33866 410576 33872
rect 409880 31204 409932 31210
rect 409880 31146 409932 31152
rect 409892 16574 409920 31146
rect 408512 16546 409184 16574
rect 409892 16546 410472 16574
rect 407212 14544 407264 14550
rect 407212 14486 407264 14492
rect 407120 3596 407172 3602
rect 407120 3538 407172 3544
rect 407224 480 407252 14486
rect 408408 3596 408460 3602
rect 408408 3538 408460 3544
rect 408420 480 408448 3538
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410444 3482 410472 16546
rect 410536 3602 410564 33866
rect 410524 3596 410576 3602
rect 410524 3538 410576 3544
rect 411904 3596 411956 3602
rect 411904 3538 411956 3544
rect 410444 3454 410840 3482
rect 410812 480 410840 3454
rect 411916 480 411944 3538
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 60007
rect 414662 57352 414718 57361
rect 414662 57287 414718 57296
rect 414296 13184 414348 13190
rect 414296 13126 414348 13132
rect 414308 480 414336 13126
rect 414676 3398 414704 57287
rect 414664 3392 414716 3398
rect 414664 3334 414716 3340
rect 415504 480 415532 77998
rect 422300 77988 422352 77994
rect 422300 77930 422352 77936
rect 418802 50280 418858 50289
rect 418802 50215 418858 50224
rect 416780 22908 416832 22914
rect 416780 22850 416832 22856
rect 416792 16574 416820 22850
rect 418160 17468 418212 17474
rect 418160 17410 418212 17416
rect 418172 16574 418200 17410
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 418816 3602 418844 50215
rect 422312 16574 422340 77930
rect 423772 69760 423824 69766
rect 423772 69702 423824 69708
rect 422942 61432 422998 61441
rect 422942 61367 422998 61376
rect 422312 16546 422616 16574
rect 420920 15904 420972 15910
rect 420920 15846 420972 15852
rect 418804 3596 418856 3602
rect 418804 3538 418856 3544
rect 420184 3596 420236 3602
rect 420184 3538 420236 3544
rect 420196 480 420224 3538
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 15846
rect 422588 480 422616 16546
rect 422956 3602 422984 61367
rect 423784 3738 423812 69702
rect 427818 43616 427874 43625
rect 427818 43551 427874 43560
rect 426440 42288 426492 42294
rect 426440 42230 426492 42236
rect 425060 25696 425112 25702
rect 425060 25638 425112 25644
rect 425072 16574 425100 25638
rect 426452 16574 426480 42230
rect 427832 16574 427860 43551
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 423772 3732 423824 3738
rect 423772 3674 423824 3680
rect 424968 3732 425020 3738
rect 424968 3674 425020 3680
rect 422944 3596 422996 3602
rect 422944 3538 422996 3544
rect 423772 3596 423824 3602
rect 423772 3538 423824 3544
rect 423784 480 423812 3538
rect 424980 480 425008 3674
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 78066
rect 432604 66904 432656 66910
rect 432604 66846 432656 66852
rect 430578 62928 430634 62937
rect 430578 62863 430634 62872
rect 430592 16574 430620 62863
rect 431960 32496 432012 32502
rect 431960 32438 432012 32444
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 3602 432000 32438
rect 432052 9104 432104 9110
rect 432052 9046 432104 9052
rect 431960 3596 432012 3602
rect 431960 3538 432012 3544
rect 432064 480 432092 9046
rect 432616 2990 432644 66846
rect 434720 29776 434772 29782
rect 434720 29718 434772 29724
rect 434732 16574 434760 29718
rect 436112 16574 436140 78639
rect 453302 75304 453358 75313
rect 453302 75239 453358 75248
rect 449900 73840 449952 73846
rect 449900 73782 449952 73788
rect 446404 72480 446456 72486
rect 446404 72422 446456 72428
rect 437478 53136 437534 53145
rect 437478 53071 437534 53080
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433248 3596 433300 3602
rect 433248 3538 433300 3544
rect 432604 2984 432656 2990
rect 432604 2926 432656 2932
rect 433260 480 433288 3538
rect 434444 2984 434496 2990
rect 434444 2926 434496 2932
rect 434456 480 434484 2926
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 53071
rect 440238 48920 440294 48929
rect 440238 48855 440294 48864
rect 439136 11824 439188 11830
rect 439136 11766 439188 11772
rect 439148 480 439176 11766
rect 440252 3602 440280 48855
rect 440332 42220 440384 42226
rect 440332 42162 440384 42168
rect 440240 3596 440292 3602
rect 440240 3538 440292 3544
rect 440344 480 440372 42162
rect 444380 40860 444432 40866
rect 444380 40802 444432 40808
rect 443000 31136 443052 31142
rect 443000 31078 443052 31084
rect 441620 17400 441672 17406
rect 441620 17342 441672 17348
rect 441632 16574 441660 17342
rect 443012 16574 443040 31078
rect 444392 16574 444420 40802
rect 445760 17332 445812 17338
rect 445760 17274 445812 17280
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 444392 16546 445064 16574
rect 441528 3596 441580 3602
rect 441528 3538 441580 3544
rect 441540 480 441568 3538
rect 442644 480 442672 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445036 480 445064 16546
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 17274
rect 446416 3602 446444 72422
rect 448520 69692 448572 69698
rect 448520 69634 448572 69640
rect 446404 3596 446456 3602
rect 446404 3538 446456 3544
rect 447416 3596 447468 3602
rect 447416 3538 447468 3544
rect 447428 480 447456 3538
rect 448532 3482 448560 69634
rect 448612 38072 448664 38078
rect 448612 38014 448664 38020
rect 448624 3602 448652 38014
rect 449912 16574 449940 73782
rect 450542 58576 450598 58585
rect 450542 58511 450598 58520
rect 449912 16546 450492 16574
rect 448612 3596 448664 3602
rect 448612 3538 448664 3544
rect 449808 3596 449860 3602
rect 449808 3538 449860 3544
rect 448532 3454 448652 3482
rect 448624 480 448652 3454
rect 449820 480 449848 3538
rect 450464 3482 450492 16546
rect 450556 4146 450584 58511
rect 450544 4140 450596 4146
rect 450544 4082 450596 4088
rect 452108 4140 452160 4146
rect 452108 4082 452160 4088
rect 450464 3454 450952 3482
rect 450924 480 450952 3454
rect 452120 480 452148 4082
rect 453316 3602 453344 75239
rect 465172 73908 465224 73914
rect 465172 73850 465224 73856
rect 459558 56128 459614 56137
rect 459558 56063 459614 56072
rect 455418 51776 455474 51785
rect 455418 51711 455474 51720
rect 454040 35352 454092 35358
rect 454040 35294 454092 35300
rect 453396 7676 453448 7682
rect 453396 7618 453448 7624
rect 453304 3596 453356 3602
rect 453304 3538 453356 3544
rect 453408 3482 453436 7618
rect 453316 3454 453436 3482
rect 453316 480 453344 3454
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454052 354 454080 35294
rect 455432 16574 455460 51711
rect 458178 46200 458234 46209
rect 458178 46135 458234 46144
rect 456892 28348 456944 28354
rect 456892 28290 456944 28296
rect 455432 16546 455736 16574
rect 455708 480 455736 16546
rect 456904 480 456932 28290
rect 458192 16574 458220 46135
rect 459572 16574 459600 56063
rect 464344 53848 464396 53854
rect 464344 53790 464396 53796
rect 463700 39500 463752 39506
rect 463700 39442 463752 39448
rect 462320 39432 462372 39438
rect 462320 39374 462372 39380
rect 460940 22840 460992 22846
rect 460940 22782 460992 22788
rect 460952 16574 460980 22782
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 458088 3528 458140 3534
rect 458088 3470 458140 3476
rect 458100 480 458128 3470
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 39374
rect 463712 16574 463740 39442
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 464356 3058 464384 53790
rect 464344 3052 464396 3058
rect 464344 2994 464396 3000
rect 465184 480 465212 73850
rect 472624 64184 472676 64190
rect 472624 64126 472676 64132
rect 466460 53100 466512 53106
rect 466460 53042 466512 53048
rect 466472 16574 466500 53042
rect 468484 51740 468536 51746
rect 468484 51682 468536 51688
rect 466472 16546 467512 16574
rect 466276 3052 466328 3058
rect 466276 2994 466328 3000
rect 466288 480 466316 2994
rect 467484 480 467512 16546
rect 468496 3534 468524 51682
rect 470598 47560 470654 47569
rect 470598 47495 470654 47504
rect 468484 3528 468536 3534
rect 468484 3470 468536 3476
rect 469864 3528 469916 3534
rect 469864 3470 469916 3476
rect 468668 3460 468720 3466
rect 468668 3402 468720 3408
rect 468680 480 468708 3402
rect 469876 480 469904 3470
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 47495
rect 471980 21480 472032 21486
rect 471980 21422 472032 21428
rect 471992 16574 472020 21422
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 472636 3534 472664 64126
rect 473452 57248 473504 57254
rect 473452 57190 473504 57196
rect 473464 16574 473492 57190
rect 474740 46300 474792 46306
rect 474740 46242 474792 46248
rect 474752 16574 474780 46242
rect 476118 43480 476174 43489
rect 476118 43415 476174 43424
rect 476132 16574 476160 43415
rect 477500 17264 477552 17270
rect 477500 17206 477552 17212
rect 477512 16574 477540 17206
rect 480272 16574 480300 78814
rect 483020 78804 483072 78810
rect 483020 78746 483072 78752
rect 480904 75404 480956 75410
rect 480904 75346 480956 75352
rect 473464 16546 474136 16574
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 477512 16546 478184 16574
rect 480272 16546 480576 16574
rect 472624 3528 472676 3534
rect 472624 3470 472676 3476
rect 473452 3528 473504 3534
rect 473452 3470 473504 3476
rect 473464 480 473492 3470
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 478156 480 478184 16546
rect 478880 15972 478932 15978
rect 478880 15914 478932 15920
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 15914
rect 480548 480 480576 16546
rect 480916 3466 480944 75346
rect 481640 38004 481692 38010
rect 481640 37946 481692 37952
rect 481652 16574 481680 37946
rect 483032 16574 483060 78746
rect 500960 78736 501012 78742
rect 500960 78678 501012 78684
rect 489182 71360 489238 71369
rect 489182 71295 489238 71304
rect 486424 54528 486476 54534
rect 486424 54470 486476 54476
rect 484400 36644 484452 36650
rect 484400 36586 484452 36592
rect 484412 16574 484440 36586
rect 481652 16546 481772 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 480904 3460 480956 3466
rect 480904 3402 480956 3408
rect 481744 480 481772 16546
rect 482836 6316 482888 6322
rect 482836 6258 482888 6264
rect 482848 480 482876 6258
rect 484044 480 484072 16546
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 486332 4888 486384 4894
rect 486332 4830 486384 4836
rect 486344 2530 486372 4830
rect 486436 3534 486464 54470
rect 488540 47660 488592 47666
rect 488540 47602 488592 47608
rect 488552 16574 488580 47602
rect 488552 16546 488856 16574
rect 486424 3528 486476 3534
rect 486424 3470 486476 3476
rect 487620 3528 487672 3534
rect 487620 3470 487672 3476
rect 486344 2502 486464 2530
rect 486436 480 486464 2502
rect 487632 480 487660 3470
rect 488828 480 488856 16546
rect 489196 4146 489224 71295
rect 498198 69728 498254 69737
rect 498198 69663 498254 69672
rect 490012 58676 490064 58682
rect 490012 58618 490064 58624
rect 490024 6914 490052 58618
rect 494058 36544 494114 36553
rect 494058 36479 494114 36488
rect 491300 33856 491352 33862
rect 491300 33798 491352 33804
rect 491312 16574 491340 33798
rect 494072 16574 494100 36479
rect 495440 31068 495492 31074
rect 495440 31010 495492 31016
rect 491312 16546 492352 16574
rect 494072 16546 494744 16574
rect 489932 6886 490052 6914
rect 489184 4140 489236 4146
rect 489184 4082 489236 4088
rect 489932 480 489960 6886
rect 491116 4140 491168 4146
rect 491116 4082 491168 4088
rect 491128 480 491156 4082
rect 492324 480 492352 16546
rect 493048 10328 493100 10334
rect 493048 10270 493100 10276
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 354 493088 10270
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 31010
rect 497096 3596 497148 3602
rect 497096 3538 497148 3544
rect 497108 480 497136 3538
rect 498212 480 498240 69663
rect 499578 55992 499634 56001
rect 499578 55927 499634 55936
rect 498292 42152 498344 42158
rect 498292 42094 498344 42100
rect 498304 16574 498332 42094
rect 499592 16574 499620 55927
rect 500972 16574 501000 78678
rect 509884 76560 509936 76566
rect 509884 76502 509936 76508
rect 506480 75336 506532 75342
rect 506480 75278 506532 75284
rect 504364 68332 504416 68338
rect 504364 68274 504416 68280
rect 502340 35284 502392 35290
rect 502340 35226 502392 35232
rect 502352 16574 502380 35226
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 503720 14476 503772 14482
rect 503720 14418 503772 14424
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 14418
rect 504376 3534 504404 68274
rect 506492 3534 506520 75278
rect 507858 71224 507914 71233
rect 507858 71159 507914 71168
rect 506572 28280 506624 28286
rect 506572 28222 506624 28228
rect 504364 3528 504416 3534
rect 504364 3470 504416 3476
rect 505376 3528 505428 3534
rect 505376 3470 505428 3476
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 505388 480 505416 3470
rect 506584 3346 506612 28222
rect 507872 16574 507900 71159
rect 509240 26988 509292 26994
rect 509240 26930 509292 26936
rect 509252 16574 509280 26930
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 509896 3534 509924 76502
rect 511264 75268 511316 75274
rect 511264 75210 511316 75216
rect 511276 16574 511304 75210
rect 514022 65648 514078 65657
rect 514022 65583 514078 65592
rect 511998 64288 512054 64297
rect 511998 64223 512054 64232
rect 511276 16546 511396 16574
rect 511264 13116 511316 13122
rect 511264 13058 511316 13064
rect 509884 3528 509936 3534
rect 509884 3470 509936 3476
rect 511276 480 511304 13058
rect 511368 3194 511396 16546
rect 511356 3188 511408 3194
rect 511356 3130 511408 3136
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 64223
rect 513380 25628 513432 25634
rect 513380 25570 513432 25576
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 25570
rect 514036 3058 514064 65583
rect 516140 40792 516192 40798
rect 516140 40734 516192 40740
rect 516152 16574 516180 40734
rect 520280 39364 520332 39370
rect 520280 39306 520332 39312
rect 518900 19984 518952 19990
rect 518900 19926 518952 19932
rect 518912 16574 518940 19926
rect 516152 16546 517192 16574
rect 518912 16546 519584 16574
rect 514760 3188 514812 3194
rect 514760 3130 514812 3136
rect 514024 3052 514076 3058
rect 514024 2994 514076 3000
rect 514772 480 514800 3130
rect 515956 3052 516008 3058
rect 515956 2994 516008 3000
rect 515968 480 515996 2994
rect 517164 480 517192 16546
rect 518348 3528 518400 3534
rect 518348 3470 518400 3476
rect 518360 480 518388 3470
rect 519556 480 519584 16546
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 39306
rect 522304 24200 522356 24206
rect 522304 24142 522356 24148
rect 521844 3460 521896 3466
rect 521844 3402 521896 3408
rect 521856 480 521884 3402
rect 522316 3126 522344 24142
rect 522396 18760 522448 18766
rect 522396 18702 522448 18708
rect 522408 3466 522436 18702
rect 523144 6914 523172 80815
rect 525798 80744 525854 80753
rect 525798 80679 525854 80688
rect 524420 26920 524472 26926
rect 524420 26862 524472 26868
rect 524432 16574 524460 26862
rect 525812 16574 525840 80679
rect 536838 78976 536894 78985
rect 536838 78911 536894 78920
rect 535458 75168 535514 75177
rect 535458 75103 535514 75112
rect 531318 71088 531374 71097
rect 531318 71023 531374 71032
rect 527822 65512 527878 65521
rect 527822 65447 527878 65456
rect 527180 44940 527232 44946
rect 527180 44882 527232 44888
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523052 6886 523172 6914
rect 522396 3460 522448 3466
rect 522396 3402 522448 3408
rect 522304 3120 522356 3126
rect 522304 3062 522356 3068
rect 523052 480 523080 6886
rect 524236 3120 524288 3126
rect 524236 3062 524288 3068
rect 524248 480 524276 3062
rect 525444 480 525472 16546
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527192 6914 527220 44882
rect 527836 16574 527864 65447
rect 529940 60852 529992 60858
rect 529940 60794 529992 60800
rect 528560 42084 528612 42090
rect 528560 42026 528612 42032
rect 527836 16546 527956 16574
rect 527192 6886 527864 6914
rect 527836 480 527864 6886
rect 527928 3534 527956 16546
rect 527916 3528 527968 3534
rect 527916 3470 527968 3476
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 42026
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 60794
rect 531332 480 531360 71023
rect 531412 25560 531464 25566
rect 531412 25502 531464 25508
rect 531424 16574 531452 25502
rect 534080 22772 534132 22778
rect 534080 22714 534132 22720
rect 534092 16574 534120 22714
rect 535472 16574 535500 75103
rect 536852 16574 536880 78911
rect 553398 76528 553454 76537
rect 553398 76463 553454 76472
rect 549260 75200 549312 75206
rect 549260 75142 549312 75148
rect 539600 66292 539652 66298
rect 539600 66234 539652 66240
rect 538220 37936 538272 37942
rect 538220 37878 538272 37884
rect 531424 16546 532096 16574
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 533712 3528 533764 3534
rect 533712 3470 533764 3476
rect 533724 480 533752 3470
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 37878
rect 539612 3534 539640 66234
rect 543738 64152 543794 64161
rect 543738 64087 543794 64096
rect 542360 44872 542412 44878
rect 542360 44814 542412 44820
rect 539692 32428 539744 32434
rect 539692 32370 539744 32376
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 32370
rect 542372 16574 542400 44814
rect 543752 16574 543780 64087
rect 547878 62792 547934 62801
rect 547878 62727 547934 62736
rect 545762 57216 545818 57225
rect 545762 57151 545818 57160
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 541992 4820 542044 4826
rect 541992 4762 542044 4768
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 4762
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 7608 545540 7614
rect 545488 7550 545540 7556
rect 545500 480 545528 7550
rect 545776 3534 545804 57151
rect 546500 24132 546552 24138
rect 546500 24074 546552 24080
rect 545764 3528 545816 3534
rect 545764 3470 545816 3476
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 24074
rect 547892 480 547920 62727
rect 549272 16574 549300 75142
rect 552020 36576 552072 36582
rect 552020 36518 552072 36524
rect 552032 16574 552060 36518
rect 553412 16574 553440 76463
rect 561678 69592 561734 69601
rect 561678 69527 561734 69536
rect 560944 67652 560996 67658
rect 560944 67594 560996 67600
rect 556160 49020 556212 49026
rect 556160 48962 556212 48968
rect 554780 29708 554832 29714
rect 554780 29650 554832 29656
rect 549272 16546 550312 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 548616 11756 548668 11762
rect 548616 11698 548668 11704
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 11698
rect 550284 480 550312 16546
rect 551468 3528 551520 3534
rect 551468 3470 551520 3476
rect 551480 480 551508 3470
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 29650
rect 556172 16574 556200 48962
rect 558184 29640 558236 29646
rect 558184 29582 558236 29588
rect 556172 16546 556936 16574
rect 556160 9036 556212 9042
rect 556160 8978 556212 8984
rect 556172 480 556200 8978
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558196 3534 558224 29582
rect 558552 6248 558604 6254
rect 558552 6190 558604 6196
rect 558184 3528 558236 3534
rect 558184 3470 558236 3476
rect 558564 480 558592 6190
rect 559748 3528 559800 3534
rect 559748 3470 559800 3476
rect 559760 480 559788 3470
rect 560956 3466 560984 67594
rect 561692 16574 561720 69527
rect 565818 68232 565874 68241
rect 565818 68167 565874 68176
rect 563702 55856 563758 55865
rect 563702 55791 563758 55800
rect 561692 16546 562088 16574
rect 560852 3460 560904 3466
rect 560852 3402 560904 3408
rect 560944 3460 560996 3466
rect 560944 3402 560996 3408
rect 560864 480 560892 3402
rect 562060 480 562088 16546
rect 563244 6180 563296 6186
rect 563244 6122 563296 6128
rect 563256 480 563284 6122
rect 563716 3534 563744 55791
rect 564532 40724 564584 40730
rect 564532 40666 564584 40672
rect 564544 6914 564572 40666
rect 565832 16574 565860 68167
rect 574744 60784 574796 60790
rect 574744 60726 574796 60732
rect 567842 59936 567898 59945
rect 567842 59871 567898 59880
rect 567200 18692 567252 18698
rect 567200 18634 567252 18640
rect 567212 16574 567240 18634
rect 565832 16546 566872 16574
rect 567212 16546 567608 16574
rect 564452 6886 564572 6914
rect 563704 3528 563756 3534
rect 563704 3470 563756 3476
rect 564452 480 564480 6886
rect 565636 3528 565688 3534
rect 565636 3470 565688 3476
rect 565648 480 565676 3470
rect 566844 480 566872 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567580 354 567608 16546
rect 567856 3534 567884 59871
rect 569960 49768 570012 49774
rect 569960 49710 570012 49716
rect 569972 16574 570000 49710
rect 571984 46232 572036 46238
rect 571984 46174 572036 46180
rect 571340 35216 571392 35222
rect 571340 35158 571392 35164
rect 569972 16546 570368 16574
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 569132 3528 569184 3534
rect 569132 3470 569184 3476
rect 569144 480 569172 3470
rect 570340 480 570368 16546
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 567998 -960 568110 326
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 35158
rect 571996 3534 572024 46174
rect 574100 18624 574152 18630
rect 574100 18566 574152 18572
rect 574112 16574 574140 18566
rect 574112 16546 574692 16574
rect 571984 3528 572036 3534
rect 571984 3470 572036 3476
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 574664 3482 574692 16546
rect 574756 3602 574784 60726
rect 576136 6866 576164 139431
rect 580276 99521 580304 146270
rect 580368 143546 580396 152623
rect 580448 146396 580500 146402
rect 580448 146338 580500 146344
rect 580356 143540 580408 143546
rect 580356 143482 580408 143488
rect 580460 139369 580488 146338
rect 580446 139360 580502 139369
rect 580446 139295 580502 139304
rect 580262 99512 580318 99521
rect 580262 99447 580318 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580998 78568 581054 78577
rect 580998 78503 581054 78512
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 578240 50380 578292 50386
rect 578240 50322 578292 50328
rect 576860 33788 576912 33794
rect 576860 33730 576912 33736
rect 576872 16574 576900 33730
rect 578252 16574 578280 50322
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 581012 16574 581040 78503
rect 582380 47592 582432 47598
rect 582380 47534 582432 47540
rect 582392 16574 582420 47534
rect 576872 16546 576992 16574
rect 578252 16546 578648 16574
rect 581012 16546 581776 16574
rect 582392 16546 583432 16574
rect 576124 6860 576176 6866
rect 576124 6802 576176 6808
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 576308 3596 576360 3602
rect 576308 3538 576360 3544
rect 572720 3460 572772 3466
rect 572720 3402 572772 3408
rect 572732 480 572760 3402
rect 573928 480 573956 3470
rect 574664 3454 575152 3482
rect 575124 480 575152 3454
rect 576320 480 576348 3538
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578620 480 578648 16546
rect 581000 8968 581052 8974
rect 581000 8910 581052 8916
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 8910
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3146 449520 3202 449576
rect 2870 410488 2926 410544
rect 2778 371340 2834 371376
rect 2778 371320 2780 371340
rect 2780 371320 2832 371340
rect 2832 371320 2834 371340
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3054 267144 3110 267200
rect 3514 462576 3570 462632
rect 3514 423544 3570 423600
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3514 358420 3570 358456
rect 3514 358400 3516 358420
rect 3516 358400 3568 358420
rect 3568 358400 3570 358420
rect 3514 306176 3570 306232
rect 3514 293120 3570 293176
rect 2778 214920 2834 214976
rect 3514 254088 3570 254144
rect 3514 241032 3570 241088
rect 3422 201864 3478 201920
rect 107382 200504 107438 200560
rect 107290 200368 107346 200424
rect 106094 199552 106150 199608
rect 102046 199008 102102 199064
rect 100574 197920 100630 197976
rect 3422 188808 3478 188864
rect 3422 162832 3478 162888
rect 3422 149776 3478 149832
rect 3146 110608 3202 110664
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3514 71612 3516 71632
rect 3516 71612 3568 71632
rect 3568 71612 3570 71632
rect 3514 71576 3570 71612
rect 3422 45464 3478 45520
rect 3422 6432 3478 6488
rect 8942 68176 8998 68232
rect 11058 66816 11114 66872
rect 31022 139440 31078 139496
rect 95238 81504 95294 81560
rect 17314 36488 17370 36544
rect 34518 76472 34574 76528
rect 25502 57160 25558 57216
rect 24858 33768 24914 33824
rect 27710 51720 27766 51776
rect 30378 50224 30434 50280
rect 41418 69536 41474 69592
rect 40038 66952 40094 67008
rect 39302 48864 39358 48920
rect 44178 47504 44234 47560
rect 57242 65456 57298 65512
rect 56598 46144 56654 46200
rect 60738 77832 60794 77888
rect 75182 62736 75238 62792
rect 74538 43424 74594 43480
rect 77298 57296 77354 57352
rect 84198 54440 84254 54496
rect 96618 75112 96674 75168
rect 100482 148280 100538 148336
rect 100758 77152 100814 77208
rect 101586 77152 101642 77208
rect 100758 76472 100814 76528
rect 100758 57840 100814 57896
rect 101678 57840 101734 57896
rect 100758 57160 100814 57216
rect 100758 52400 100814 52456
rect 100758 51720 100814 51776
rect 100850 50904 100906 50960
rect 100850 50224 100906 50280
rect 101862 50904 101918 50960
rect 100850 49544 100906 49600
rect 101770 49544 101826 49600
rect 100850 48864 100906 48920
rect 104254 196968 104310 197024
rect 102874 69536 102930 69592
rect 102046 52400 102102 52456
rect 100850 48184 100906 48240
rect 101954 48184 102010 48240
rect 100850 47504 100906 47560
rect 104714 193840 104770 193896
rect 104254 67496 104310 67552
rect 105450 66136 105506 66192
rect 105450 65456 105506 65512
rect 105726 80144 105782 80200
rect 105634 72936 105690 72992
rect 107566 198736 107622 198792
rect 107474 196832 107530 196888
rect 106738 75656 106794 75712
rect 108302 192480 108358 192536
rect 106186 66136 106242 66192
rect 108394 44104 108450 44160
rect 108394 43424 108450 43480
rect 110970 189624 111026 189680
rect 110418 63416 110474 63472
rect 110418 62736 110474 62792
rect 110326 57296 110382 57352
rect 111338 192616 111394 192672
rect 110970 75520 111026 75576
rect 112350 192752 112406 192808
rect 111706 63416 111762 63472
rect 112534 74024 112590 74080
rect 111798 55120 111854 55176
rect 113086 55120 113142 55176
rect 111798 54440 111854 54496
rect 110510 46824 110566 46880
rect 110878 46824 110934 46880
rect 110510 46144 110566 46200
rect 113730 138896 113786 138952
rect 113730 76608 113786 76664
rect 114282 195336 114338 195392
rect 114466 71304 114522 71360
rect 114374 68856 114430 68912
rect 114926 73888 114982 73944
rect 114834 68720 114890 68776
rect 115110 139032 115166 139088
rect 115110 69944 115166 70000
rect 115662 77016 115718 77072
rect 116306 144608 116362 144664
rect 115754 74976 115810 75032
rect 116398 80688 116454 80744
rect 116306 71712 116362 71768
rect 117042 76880 117098 76936
rect 117134 72664 117190 72720
rect 116766 71440 116822 71496
rect 111614 3304 111670 3360
rect 117962 146920 118018 146976
rect 118422 146920 118478 146976
rect 118330 144744 118386 144800
rect 117962 79464 118018 79520
rect 118606 196696 118662 196752
rect 118606 72800 118662 72856
rect 119342 142704 119398 142760
rect 119986 200640 120042 200696
rect 119618 138624 119674 138680
rect 119526 75792 119582 75848
rect 129830 262248 129886 262304
rect 132038 261024 132094 261080
rect 135902 265104 135958 265160
rect 137466 260888 137522 260944
rect 138754 264968 138810 265024
rect 138662 262792 138718 262848
rect 140318 262656 140374 262712
rect 139674 260344 139730 260400
rect 140778 260072 140834 260128
rect 141744 260072 141800 260128
rect 142434 260072 142490 260128
rect 143630 260208 143686 260264
rect 143400 260072 143456 260128
rect 144504 260208 144560 260264
rect 146206 263880 146262 263936
rect 145286 263608 145342 263664
rect 145562 263608 145618 263664
rect 147770 263744 147826 263800
rect 146942 262520 146998 262576
rect 148506 262928 148562 262984
rect 144918 259800 144974 259856
rect 146482 259664 146538 259720
rect 150530 262384 150586 262440
rect 153382 275984 153438 276040
rect 156050 277480 156106 277536
rect 157338 260208 157394 260264
rect 158810 262656 158866 262712
rect 158304 260208 158360 260264
rect 159914 262656 159970 262712
rect 160098 259936 160154 259992
rect 162214 265512 162270 265568
rect 162030 262384 162086 262440
rect 161478 260752 161534 260808
rect 160926 259936 160982 259992
rect 163502 265104 163558 265160
rect 163410 263200 163466 263256
rect 163410 262520 163466 262576
rect 162674 260752 162730 260808
rect 162582 259800 162638 259856
rect 163594 263200 163650 263256
rect 164882 264968 164938 265024
rect 165158 265240 165214 265296
rect 165158 264968 165214 265024
rect 167458 265512 167514 265568
rect 167550 265376 167606 265432
rect 167458 265104 167514 265160
rect 158626 259664 158682 259720
rect 149058 259528 149114 259584
rect 149794 259528 149850 259584
rect 155222 259528 155278 259584
rect 185674 259528 185730 259584
rect 120814 142160 120870 142216
rect 121090 76744 121146 76800
rect 121918 147736 121974 147792
rect 121642 85176 121698 85232
rect 121182 75384 121238 75440
rect 122194 128424 122250 128480
rect 122194 123120 122250 123176
rect 121918 122712 121974 122768
rect 121918 113328 121974 113384
rect 122102 122712 122158 122768
rect 122194 122440 122250 122496
rect 122194 113464 122250 113520
rect 122102 113192 122158 113248
rect 122194 112784 122250 112840
rect 122194 103808 122250 103864
rect 121918 103264 121974 103320
rect 121918 94016 121974 94072
rect 122102 103400 122158 103456
rect 122194 103128 122250 103184
rect 122194 94152 122250 94208
rect 122102 93880 122158 93936
rect 122010 85176 122066 85232
rect 121918 75112 121974 75168
rect 122194 93472 122250 93528
rect 122194 89664 122250 89720
rect 122378 85040 122434 85096
rect 122378 84632 122434 84688
rect 122470 80280 122526 80336
rect 122654 75248 122710 75304
rect 122470 74568 122526 74624
rect 123850 199280 123906 199336
rect 123758 199144 123814 199200
rect 123206 139576 123262 139632
rect 123298 138760 123354 138816
rect 123482 140256 123538 140312
rect 123850 72528 123906 72584
rect 127622 200232 127678 200288
rect 124034 142160 124090 142216
rect 124954 148416 125010 148472
rect 126702 197376 126758 197432
rect 125506 140800 125562 140856
rect 126242 140936 126298 140992
rect 125046 139576 125102 139632
rect 126610 140256 126666 140312
rect 124954 139304 125010 139360
rect 126150 139340 126152 139360
rect 126152 139340 126204 139360
rect 126204 139340 126206 139360
rect 126150 139304 126206 139340
rect 128082 193840 128138 193896
rect 127622 140120 127678 140176
rect 129002 199824 129058 199880
rect 129002 196424 129058 196480
rect 128726 195336 128782 195392
rect 130474 200404 130476 200424
rect 130476 200404 130528 200424
rect 130528 200404 130530 200424
rect 130474 200368 130530 200404
rect 131302 200368 131358 200424
rect 130014 200096 130070 200152
rect 131302 200096 131358 200152
rect 129554 199552 129610 199608
rect 129278 199008 129334 199064
rect 132038 200640 132094 200696
rect 132222 200660 132278 200696
rect 132222 200640 132224 200660
rect 132224 200640 132276 200660
rect 132276 200640 132278 200660
rect 178682 200640 178738 200696
rect 131670 200096 131726 200152
rect 131762 199824 131818 199880
rect 131578 199688 131634 199744
rect 130290 146240 130346 146296
rect 129830 146104 129886 146160
rect 129738 145968 129794 146024
rect 130474 197104 130530 197160
rect 132222 199980 132278 200016
rect 132222 199960 132224 199980
rect 132224 199960 132276 199980
rect 132276 199960 132278 199980
rect 132130 199844 132186 199880
rect 132130 199824 132132 199844
rect 132132 199824 132184 199844
rect 132184 199824 132186 199844
rect 132912 199824 132968 199880
rect 132498 199552 132554 199608
rect 132682 196152 132738 196208
rect 133372 199824 133428 199880
rect 132406 196016 132462 196072
rect 132866 196016 132922 196072
rect 133326 197784 133382 197840
rect 133326 197648 133382 197704
rect 133648 199824 133704 199880
rect 133924 199824 133980 199880
rect 133510 198600 133566 198656
rect 133694 197920 133750 197976
rect 133878 197784 133934 197840
rect 134430 199688 134486 199744
rect 134430 197920 134486 197976
rect 134522 196968 134578 197024
rect 132682 148280 132738 148336
rect 132590 143248 132646 143304
rect 135488 199824 135544 199880
rect 135442 199688 135498 199744
rect 135258 198464 135314 198520
rect 135166 197920 135222 197976
rect 135258 197376 135314 197432
rect 135534 199008 135590 199064
rect 135718 191120 135774 191176
rect 136500 199824 136556 199880
rect 136546 199688 136602 199744
rect 136776 199824 136832 199880
rect 137052 199824 137108 199880
rect 136454 199552 136510 199608
rect 136638 199588 136640 199608
rect 136640 199588 136692 199608
rect 136692 199588 136694 199608
rect 136638 199552 136694 199588
rect 136454 199008 136510 199064
rect 136546 198736 136602 198792
rect 136546 198056 136602 198112
rect 136822 199688 136878 199744
rect 135994 190984 136050 191040
rect 137696 199824 137752 199880
rect 137880 199824 137936 199880
rect 138064 199824 138120 199880
rect 138248 199824 138304 199880
rect 138432 199824 138488 199880
rect 138984 199824 139040 199880
rect 137374 197920 137430 197976
rect 137098 195064 137154 195120
rect 137650 197784 137706 197840
rect 138110 199552 138166 199608
rect 138294 199552 138350 199608
rect 138570 196832 138626 196888
rect 137282 149640 137338 149696
rect 138938 199688 138994 199744
rect 139444 199858 139500 199914
rect 140088 199824 140144 199880
rect 139490 199552 139546 199608
rect 139306 199008 139362 199064
rect 139490 198736 139546 198792
rect 139398 198056 139454 198112
rect 139950 198600 140006 198656
rect 139858 198056 139914 198112
rect 140272 199708 140328 199710
rect 140272 199656 140274 199708
rect 140274 199656 140326 199708
rect 140326 199656 140328 199708
rect 140272 199654 140328 199656
rect 140318 198056 140374 198112
rect 140824 199688 140880 199744
rect 141008 199824 141064 199880
rect 141284 199824 141340 199880
rect 141560 199824 141616 199880
rect 140686 199008 140742 199064
rect 138754 183232 138810 183288
rect 141514 199688 141570 199744
rect 141330 199552 141386 199608
rect 141330 192616 141386 192672
rect 140870 144472 140926 144528
rect 138662 143928 138718 143984
rect 139398 143792 139454 143848
rect 140318 141752 140374 141808
rect 142112 199858 142168 199914
rect 141606 192752 141662 192808
rect 142480 199858 142536 199914
rect 141974 196016 142030 196072
rect 141974 195336 142030 195392
rect 141974 195064 142030 195120
rect 142710 199552 142766 199608
rect 141790 188808 141846 188864
rect 143170 199688 143226 199744
rect 143492 199824 143548 199880
rect 142802 192480 142858 192536
rect 143446 199008 143502 199064
rect 144504 199858 144560 199914
rect 143814 197512 143870 197568
rect 143538 194112 143594 194168
rect 144090 198872 144146 198928
rect 144182 198736 144238 198792
rect 144090 195336 144146 195392
rect 143998 193160 144054 193216
rect 144366 198464 144422 198520
rect 145424 199858 145480 199914
rect 146160 199824 146216 199880
rect 144918 197920 144974 197976
rect 145378 198328 145434 198384
rect 145562 197784 145618 197840
rect 141514 141208 141570 141264
rect 141422 141072 141478 141128
rect 142250 141616 142306 141672
rect 143630 141480 143686 141536
rect 145010 143112 145066 143168
rect 146114 195472 146170 195528
rect 145654 148416 145710 148472
rect 146758 197920 146814 197976
rect 146482 197240 146538 197296
rect 146666 145832 146722 145888
rect 146298 145696 146354 145752
rect 145838 144336 145894 144392
rect 146390 142840 146446 142896
rect 147540 199858 147596 199914
rect 147816 199824 147872 199880
rect 148000 199858 148056 199914
rect 148184 199858 148240 199914
rect 147034 199008 147090 199064
rect 147218 198872 147274 198928
rect 147218 198736 147274 198792
rect 146850 195744 146906 195800
rect 148414 199688 148470 199744
rect 148552 199724 148554 199744
rect 148554 199724 148606 199744
rect 148606 199724 148608 199744
rect 148552 199688 148608 199724
rect 147678 199552 147734 199608
rect 147954 198892 148010 198928
rect 147954 198872 147956 198892
rect 147956 198872 148008 198892
rect 148008 198872 148010 198892
rect 148138 198872 148194 198928
rect 148736 199688 148792 199744
rect 148414 199552 148470 199608
rect 147586 147056 147642 147112
rect 148782 199588 148784 199608
rect 148784 199588 148836 199608
rect 148836 199588 148838 199608
rect 148782 199552 148838 199588
rect 148598 191120 148654 191176
rect 147678 145560 147734 145616
rect 148046 142976 148102 143032
rect 149380 199858 149436 199914
rect 149656 199858 149712 199914
rect 149932 199824 149988 199880
rect 148966 199452 148968 199472
rect 148968 199452 149020 199472
rect 149020 199452 149022 199472
rect 148966 199416 149022 199452
rect 149058 190984 149114 191040
rect 149426 198464 149482 198520
rect 149610 199416 149666 199472
rect 149518 193976 149574 194032
rect 149886 199144 149942 199200
rect 150760 199858 150816 199914
rect 151220 199824 151276 199880
rect 151404 199824 151460 199880
rect 150070 196968 150126 197024
rect 149794 196424 149850 196480
rect 150438 199280 150494 199336
rect 150346 195608 150402 195664
rect 150806 195608 150862 195664
rect 149702 142704 149758 142760
rect 150622 146920 150678 146976
rect 150438 141344 150494 141400
rect 151266 196016 151322 196072
rect 152048 199824 152104 199880
rect 151726 199416 151782 199472
rect 152002 197104 152058 197160
rect 152508 199858 152564 199914
rect 152784 199858 152840 199914
rect 153060 199858 153116 199914
rect 153612 199824 153668 199880
rect 152646 196560 152702 196616
rect 152186 183504 152242 183560
rect 151726 149640 151782 149696
rect 150990 144064 151046 144120
rect 154164 199824 154220 199880
rect 154440 199824 154496 199880
rect 152554 144200 152610 144256
rect 153658 197376 153714 197432
rect 153658 190848 153714 190904
rect 154026 199280 154082 199336
rect 154026 191256 154082 191312
rect 153842 189352 153898 189408
rect 154808 199824 154864 199880
rect 155268 199858 155324 199914
rect 154854 199452 154856 199472
rect 154856 199452 154908 199472
rect 154908 199452 154910 199472
rect 154854 199416 154910 199452
rect 154578 198600 154634 198656
rect 154578 198328 154634 198384
rect 154946 199280 155002 199336
rect 154946 198600 155002 198656
rect 154854 195336 154910 195392
rect 155038 193976 155094 194032
rect 155820 199824 155876 199880
rect 153658 142160 153714 142216
rect 155774 199280 155830 199336
rect 155038 150048 155094 150104
rect 154854 149776 154910 149832
rect 155314 142704 155370 142760
rect 154762 139984 154818 140040
rect 157016 199858 157072 199914
rect 156510 198056 156566 198112
rect 156970 199416 157026 199472
rect 156878 198872 156934 198928
rect 156970 198736 157026 198792
rect 157154 199280 157210 199336
rect 156418 144200 156474 144256
rect 156970 142840 157026 142896
rect 156510 140120 156566 140176
rect 157430 198192 157486 198248
rect 157430 197648 157486 197704
rect 157522 196832 157578 196888
rect 157338 195200 157394 195256
rect 157890 198736 157946 198792
rect 157706 196696 157762 196752
rect 158258 199144 158314 199200
rect 158258 198192 158314 198248
rect 157154 149912 157210 149968
rect 157430 147328 157486 147384
rect 158534 199280 158590 199336
rect 158534 199144 158590 199200
rect 158902 199416 158958 199472
rect 160236 199824 160292 199880
rect 158810 195608 158866 195664
rect 158534 150184 158590 150240
rect 159178 197512 159234 197568
rect 159454 196560 159510 196616
rect 159730 196696 159786 196752
rect 158074 145696 158130 145752
rect 158074 144064 158130 144120
rect 160190 195472 160246 195528
rect 161018 197240 161074 197296
rect 161294 197376 161350 197432
rect 161892 199824 161948 199880
rect 160742 190440 160798 190496
rect 161386 190304 161442 190360
rect 161386 180784 161442 180840
rect 161386 180648 161442 180704
rect 161386 171128 161442 171184
rect 161386 170992 161442 171048
rect 161386 161472 161442 161528
rect 161386 161336 161442 161392
rect 161386 151816 161442 151872
rect 161386 151680 161442 151736
rect 160558 144336 160614 144392
rect 160006 142976 160062 143032
rect 161662 198328 161718 198384
rect 162628 199824 162684 199880
rect 163456 199824 163512 199880
rect 163824 199824 163880 199880
rect 162122 199280 162178 199336
rect 162490 196696 162546 196752
rect 163042 197512 163098 197568
rect 161662 152360 161718 152416
rect 162766 144472 162822 144528
rect 161938 143248 161994 143304
rect 161386 142296 161442 142352
rect 161478 142024 161534 142080
rect 162950 191120 163006 191176
rect 163134 152496 163190 152552
rect 163410 197376 163466 197432
rect 163594 189352 163650 189408
rect 164238 197240 164294 197296
rect 164836 199824 164892 199880
rect 165112 199824 165168 199880
rect 164238 191120 164294 191176
rect 164882 197240 164938 197296
rect 165388 199824 165444 199880
rect 165158 199280 165214 199336
rect 165066 197512 165122 197568
rect 164974 196832 165030 196888
rect 165250 197376 165306 197432
rect 165342 197240 165398 197296
rect 164698 191120 164754 191176
rect 164606 152632 164662 152688
rect 165986 199008 166042 199064
rect 165986 198892 166042 198928
rect 165986 198872 165988 198892
rect 165988 198872 166040 198892
rect 166040 198872 166042 198892
rect 166400 199824 166456 199880
rect 166768 199824 166824 199880
rect 166354 199280 166410 199336
rect 166354 197240 166410 197296
rect 167136 199824 167192 199880
rect 167412 199824 167468 199880
rect 166814 198872 166870 198928
rect 166538 198056 166594 198112
rect 166906 196696 166962 196752
rect 167872 199824 167928 199880
rect 167550 197512 167606 197568
rect 167826 198872 167882 198928
rect 168010 197376 168066 197432
rect 167918 193840 167974 193896
rect 168286 197240 168342 197296
rect 168194 197104 168250 197160
rect 168562 193976 168618 194032
rect 169022 197376 169078 197432
rect 169298 197920 169354 197976
rect 169620 199824 169676 199880
rect 170448 199824 170504 199880
rect 169574 197240 169630 197296
rect 170402 199280 170458 199336
rect 170402 197240 170458 197296
rect 164238 145560 164294 145616
rect 163962 143928 164018 143984
rect 163594 143112 163650 143168
rect 162858 141344 162914 141400
rect 168010 144744 168066 144800
rect 166354 144608 166410 144664
rect 165250 143384 165306 143440
rect 171092 199824 171148 199880
rect 170862 199280 170918 199336
rect 170678 197376 170734 197432
rect 171552 199824 171608 199880
rect 171920 199824 171976 199880
rect 171138 199280 171194 199336
rect 171046 198192 171102 198248
rect 170034 140256 170090 140312
rect 171782 197376 171838 197432
rect 172150 199280 172206 199336
rect 172058 199008 172114 199064
rect 172472 199824 172528 199880
rect 172334 197376 172390 197432
rect 172794 199280 172850 199336
rect 172702 199008 172758 199064
rect 172702 198600 172758 198656
rect 171230 140120 171286 140176
rect 172702 147192 172758 147248
rect 172978 199280 173034 199336
rect 172886 197784 172942 197840
rect 172978 197240 173034 197296
rect 173760 199824 173816 199880
rect 173254 198772 173256 198792
rect 173256 198772 173308 198792
rect 173308 198772 173310 198792
rect 173254 198736 173310 198772
rect 173162 197240 173218 197296
rect 173162 192616 173218 192672
rect 173438 198464 173494 198520
rect 173530 197376 173586 197432
rect 174220 199824 174276 199880
rect 173714 197920 173770 197976
rect 174266 199416 174322 199472
rect 174174 198736 174230 198792
rect 174450 199008 174506 199064
rect 174358 197512 174414 197568
rect 175048 199824 175104 199880
rect 175600 199824 175656 199880
rect 174358 192480 174414 192536
rect 174818 199416 174874 199472
rect 174818 198328 174874 198384
rect 175002 197920 175058 197976
rect 174910 197376 174966 197432
rect 175002 197240 175058 197296
rect 175094 195744 175150 195800
rect 175186 195200 175242 195256
rect 174174 147600 174230 147656
rect 174358 147464 174414 147520
rect 174082 146104 174138 146160
rect 175462 199008 175518 199064
rect 175462 197240 175518 197296
rect 176014 197376 176070 197432
rect 175370 145968 175426 146024
rect 176612 199824 176668 199880
rect 176796 199824 176852 199880
rect 176198 199008 176254 199064
rect 176290 195608 176346 195664
rect 176474 199008 176530 199064
rect 176566 198464 176622 198520
rect 176750 197104 176806 197160
rect 176842 195880 176898 195936
rect 176566 192752 176622 192808
rect 175554 145832 175610 145888
rect 176658 141208 176714 141264
rect 177302 199280 177358 199336
rect 177394 198056 177450 198112
rect 177486 197920 177542 197976
rect 178314 200096 178370 200152
rect 177854 199824 177910 199880
rect 177118 195064 177174 195120
rect 178130 198464 178186 198520
rect 177762 193024 177818 193080
rect 177026 192888 177082 192944
rect 176750 141072 176806 141128
rect 178222 142160 178278 142216
rect 178038 140120 178094 140176
rect 171230 139712 171286 139768
rect 179694 193160 179750 193216
rect 179142 150320 179198 150376
rect 179142 139984 179198 140040
rect 180154 141480 180210 141536
rect 180798 140664 180854 140720
rect 181166 140664 181222 140720
rect 181810 139848 181866 139904
rect 181902 139712 181958 139768
rect 181902 139576 181958 139632
rect 181258 139440 181314 139496
rect 182822 139440 182878 139496
rect 183834 144880 183890 144936
rect 183926 140664 183982 140720
rect 184386 140392 184442 140448
rect 185030 143248 185086 143304
rect 185030 142704 185086 142760
rect 184754 140664 184810 140720
rect 185950 143384 186006 143440
rect 185858 140528 185914 140584
rect 185766 139712 185822 139768
rect 184662 139440 184718 139496
rect 126702 139304 126758 139360
rect 128266 139304 128322 139360
rect 132222 139304 132278 139360
rect 133050 139304 133106 139360
rect 145746 139304 145802 139360
rect 150898 139304 150954 139360
rect 154026 139304 154082 139360
rect 155682 139304 155738 139360
rect 155866 139304 155922 139360
rect 157062 139304 157118 139360
rect 159546 139304 159602 139360
rect 159730 139304 159786 139360
rect 178406 139304 178462 139360
rect 178866 139304 178922 139360
rect 180246 139304 180302 139360
rect 179326 80688 179382 80744
rect 179602 80688 179658 80744
rect 179878 80688 179934 80744
rect 124126 79328 124182 79384
rect 130934 80280 130990 80336
rect 130198 79872 130254 79928
rect 130106 79328 130162 79384
rect 130014 78104 130070 78160
rect 129738 75792 129794 75848
rect 128910 70080 128966 70136
rect 130382 76472 130438 76528
rect 130290 76336 130346 76392
rect 130382 75928 130438 75984
rect 130842 78532 130898 78568
rect 130842 78512 130844 78532
rect 130844 78512 130896 78532
rect 130896 78512 130898 78532
rect 131026 75792 131082 75848
rect 131946 80552 132002 80608
rect 177762 80552 177818 80608
rect 131854 80008 131910 80064
rect 178130 80416 178186 80472
rect 132222 79736 132278 79792
rect 132544 79906 132600 79962
rect 132728 79872 132784 79928
rect 133004 79906 133060 79962
rect 132682 79736 132738 79792
rect 132130 79600 132186 79656
rect 131670 75928 131726 75984
rect 132590 78104 132646 78160
rect 133326 79736 133382 79792
rect 132866 78512 132922 78568
rect 133050 78512 133106 78568
rect 132222 68176 132278 68232
rect 132958 78376 133014 78432
rect 132958 78104 133014 78160
rect 133924 79908 133926 79928
rect 133926 79908 133978 79928
rect 133978 79908 133980 79928
rect 133924 79872 133980 79908
rect 134844 79872 134900 79928
rect 135028 79906 135084 79962
rect 135396 79906 135452 79962
rect 133510 76608 133566 76664
rect 133602 76472 133658 76528
rect 134522 79736 134578 79792
rect 134062 77444 134118 77480
rect 134062 77424 134064 77444
rect 134064 77424 134116 77444
rect 134116 77424 134118 77444
rect 134062 76336 134118 76392
rect 134246 76608 134302 76664
rect 134154 74160 134210 74216
rect 134522 77152 134578 77208
rect 135120 79770 135176 79826
rect 135258 79736 135314 79792
rect 135074 79600 135130 79656
rect 134706 75928 134762 75984
rect 136408 79906 136464 79962
rect 135718 79636 135720 79656
rect 135720 79636 135772 79656
rect 135772 79636 135774 79656
rect 135718 79600 135774 79636
rect 135442 75928 135498 75984
rect 135350 75792 135406 75848
rect 135626 78512 135682 78568
rect 135810 77832 135866 77888
rect 135994 78240 136050 78296
rect 135902 75928 135958 75984
rect 136776 79906 136832 79962
rect 136362 79600 136418 79656
rect 137052 79906 137108 79962
rect 136914 77696 136970 77752
rect 137098 79756 137154 79792
rect 137328 79872 137384 79928
rect 137098 79736 137100 79756
rect 137100 79736 137152 79756
rect 137152 79736 137154 79756
rect 136730 74840 136786 74896
rect 137282 78240 137338 78296
rect 137880 79872 137936 79928
rect 138340 79906 138396 79962
rect 137650 79600 137706 79656
rect 137558 77288 137614 77344
rect 137926 78512 137982 78568
rect 138294 79736 138350 79792
rect 138708 79872 138764 79928
rect 138110 78512 138166 78568
rect 138294 78648 138350 78704
rect 138018 77696 138074 77752
rect 138202 77832 138258 77888
rect 138110 77444 138166 77480
rect 138110 77424 138112 77444
rect 138112 77424 138164 77444
rect 138164 77424 138166 77444
rect 138294 77424 138350 77480
rect 138202 77288 138258 77344
rect 139352 79906 139408 79962
rect 139030 79600 139086 79656
rect 138754 77560 138810 77616
rect 139536 79872 139592 79928
rect 139812 79872 139868 79928
rect 139214 79636 139216 79656
rect 139216 79636 139268 79656
rect 139268 79636 139270 79656
rect 139214 79600 139270 79636
rect 139306 78104 139362 78160
rect 139306 77560 139362 77616
rect 139674 79600 139730 79656
rect 140088 79838 140144 79894
rect 139582 78920 139638 78976
rect 139674 78648 139730 78704
rect 139582 77288 139638 77344
rect 139766 77696 139822 77752
rect 140640 79872 140696 79928
rect 140824 79872 140880 79928
rect 140778 79600 140834 79656
rect 140686 78920 140742 78976
rect 140870 78920 140926 78976
rect 141192 79736 141248 79792
rect 140870 77424 140926 77480
rect 141744 79872 141800 79928
rect 141422 79620 141478 79656
rect 141422 79600 141424 79620
rect 141424 79600 141476 79620
rect 141476 79600 141478 79620
rect 141330 77152 141386 77208
rect 141928 79736 141984 79792
rect 142480 79906 142536 79962
rect 141698 79600 141754 79656
rect 142204 79736 142260 79792
rect 142526 79736 142582 79792
rect 142848 79838 142904 79894
rect 142434 79600 142490 79656
rect 141974 77424 142030 77480
rect 142066 70352 142122 70408
rect 142618 79600 142674 79656
rect 142618 77152 142674 77208
rect 142066 64912 142122 64968
rect 142066 64776 142122 64832
rect 142066 55256 142122 55312
rect 142066 55120 142122 55176
rect 142066 45600 142122 45656
rect 142066 45464 142122 45520
rect 143308 79872 143364 79928
rect 143492 79872 143548 79928
rect 142066 35944 142122 36000
rect 142066 35808 142122 35864
rect 142066 26288 142122 26344
rect 142066 26152 142122 26208
rect 142066 16632 142122 16688
rect 142066 16496 142122 16552
rect 142066 6976 142122 7032
rect 142066 6840 142122 6896
rect 143768 79872 143824 79928
rect 144780 79906 144836 79962
rect 143538 79600 143594 79656
rect 143814 78920 143870 78976
rect 143722 78648 143778 78704
rect 144688 79736 144744 79792
rect 145240 79906 145296 79962
rect 145608 79872 145664 79928
rect 145976 79872 146032 79928
rect 146160 79872 146216 79928
rect 146620 79872 146676 79928
rect 144366 79600 144422 79656
rect 144550 74704 144606 74760
rect 144826 79192 144882 79248
rect 144734 75112 144790 75168
rect 144734 71032 144790 71088
rect 145746 79756 145802 79792
rect 145746 79736 145748 79756
rect 145748 79736 145800 79756
rect 145800 79736 145802 79756
rect 145930 79736 145986 79792
rect 146114 79736 146170 79792
rect 146896 79906 146952 79962
rect 147264 79872 147320 79928
rect 145930 75384 145986 75440
rect 146114 75248 146170 75304
rect 145838 73888 145894 73944
rect 146482 79600 146538 79656
rect 146942 79736 146998 79792
rect 146758 78512 146814 78568
rect 146942 77560 146998 77616
rect 142066 3304 142122 3360
rect 147126 79192 147182 79248
rect 147586 79600 147642 79656
rect 147310 76880 147366 76936
rect 147218 69944 147274 70000
rect 147494 79056 147550 79112
rect 148460 79906 148516 79962
rect 148644 79906 148700 79962
rect 148920 79872 148976 79928
rect 148046 79756 148102 79792
rect 148046 79736 148048 79756
rect 148048 79736 148100 79756
rect 148100 79736 148102 79756
rect 148230 79736 148286 79792
rect 147678 77016 147734 77072
rect 148414 77696 148470 77752
rect 148138 75928 148194 75984
rect 148322 68856 148378 68912
rect 149104 79872 149160 79928
rect 148782 78240 148838 78296
rect 149242 79600 149298 79656
rect 148966 79056 149022 79112
rect 149150 79056 149206 79112
rect 150208 79872 150264 79928
rect 150392 79872 150448 79928
rect 149426 77832 149482 77888
rect 149702 79600 149758 79656
rect 150254 79772 150256 79792
rect 150256 79772 150308 79792
rect 150308 79772 150310 79792
rect 150254 79736 150310 79772
rect 150852 79906 150908 79962
rect 151128 79892 151184 79928
rect 151128 79872 151130 79892
rect 151130 79872 151182 79892
rect 151182 79872 151184 79892
rect 150898 79736 150954 79792
rect 151036 79736 151092 79792
rect 150162 78240 150218 78296
rect 150070 78104 150126 78160
rect 149794 50632 149850 50688
rect 150530 79620 150586 79656
rect 150530 79600 150532 79620
rect 150532 79600 150584 79620
rect 150584 79600 150586 79620
rect 150806 79328 150862 79384
rect 151082 79600 151138 79656
rect 151680 79906 151736 79962
rect 151864 79906 151920 79962
rect 151266 79620 151322 79656
rect 151266 79600 151268 79620
rect 151268 79600 151320 79620
rect 151320 79600 151322 79620
rect 151174 78648 151230 78704
rect 151450 79328 151506 79384
rect 151450 78104 151506 78160
rect 151910 79600 151966 79656
rect 151726 78376 151782 78432
rect 151634 76336 151690 76392
rect 152232 79736 152288 79792
rect 152508 79838 152564 79894
rect 152186 79348 152242 79384
rect 152186 79328 152188 79348
rect 152188 79328 152240 79348
rect 152240 79328 152242 79348
rect 152370 78512 152426 78568
rect 152278 74432 152334 74488
rect 152278 73616 152334 73672
rect 152646 79600 152702 79656
rect 152738 79464 152794 79520
rect 153014 78240 153070 78296
rect 152922 77832 152978 77888
rect 152830 76200 152886 76256
rect 152738 73616 152794 73672
rect 153106 78104 153162 78160
rect 153106 77560 153162 77616
rect 153888 79872 153944 79928
rect 153750 79600 153806 79656
rect 153474 79464 153530 79520
rect 154440 79872 154496 79928
rect 154210 79600 154266 79656
rect 154302 79464 154358 79520
rect 154210 79328 154266 79384
rect 154026 78512 154082 78568
rect 154118 77832 154174 77888
rect 153934 76608 153990 76664
rect 154578 79736 154634 79792
rect 154486 78512 154542 78568
rect 154992 79872 155048 79928
rect 154578 76880 154634 76936
rect 154578 68176 154634 68232
rect 155222 79772 155270 79792
rect 155270 79772 155278 79792
rect 155222 79736 155278 79772
rect 155544 79872 155600 79928
rect 155820 79872 155876 79928
rect 155130 78512 155186 78568
rect 155406 77832 155462 77888
rect 155590 79600 155646 79656
rect 155314 74976 155370 75032
rect 155314 73752 155370 73808
rect 155774 79464 155830 79520
rect 155682 74160 155738 74216
rect 155958 72936 156014 72992
rect 156372 79736 156428 79792
rect 156648 79736 156704 79792
rect 157016 79872 157072 79928
rect 156326 78104 156382 78160
rect 156326 77560 156382 77616
rect 156326 73072 156382 73128
rect 156050 70216 156106 70272
rect 156050 69808 156106 69864
rect 156510 77832 156566 77888
rect 157200 79872 157256 79928
rect 156786 78376 156842 78432
rect 156970 79600 157026 79656
rect 156970 78648 157026 78704
rect 156602 72256 156658 72312
rect 157062 76744 157118 76800
rect 156878 71712 156934 71768
rect 156786 69808 156842 69864
rect 157154 72936 157210 72992
rect 157752 79872 157808 79928
rect 157706 79736 157762 79792
rect 157430 77696 157486 77752
rect 157430 75248 157486 75304
rect 158580 79872 158636 79928
rect 157798 79600 157854 79656
rect 157798 79484 157854 79520
rect 157798 79464 157800 79484
rect 157800 79464 157852 79484
rect 157852 79464 157854 79484
rect 157430 72392 157486 72448
rect 158074 79636 158076 79656
rect 158076 79636 158128 79656
rect 158128 79636 158130 79656
rect 158074 79600 158130 79636
rect 158166 78648 158222 78704
rect 157982 74296 158038 74352
rect 158856 79736 158912 79792
rect 158258 74296 158314 74352
rect 158074 74024 158130 74080
rect 158534 78648 158590 78704
rect 158718 79192 158774 79248
rect 158626 77832 158682 77888
rect 158626 74024 158682 74080
rect 158626 73752 158682 73808
rect 159086 79192 159142 79248
rect 159500 79906 159556 79962
rect 159684 79872 159740 79928
rect 159408 79736 159464 79792
rect 159960 79906 160016 79962
rect 159638 79600 159694 79656
rect 159822 71712 159878 71768
rect 160328 79872 160384 79928
rect 160236 79736 160292 79792
rect 160190 79056 160246 79112
rect 160006 78376 160062 78432
rect 158718 21256 158774 21312
rect 160742 79756 160798 79792
rect 160742 79736 160744 79756
rect 160744 79736 160796 79756
rect 160796 79736 160798 79756
rect 161432 79872 161488 79928
rect 160558 79056 160614 79112
rect 160466 78648 160522 78704
rect 160558 77968 160614 78024
rect 160926 79620 160982 79656
rect 160926 79600 160928 79620
rect 160928 79600 160980 79620
rect 160980 79600 160982 79620
rect 160834 77288 160890 77344
rect 161202 79736 161258 79792
rect 161708 79872 161764 79928
rect 161110 77288 161166 77344
rect 160098 15816 160154 15872
rect 161662 78784 161718 78840
rect 162444 79872 162500 79928
rect 162720 79872 162776 79928
rect 162904 79906 162960 79962
rect 161846 79056 161902 79112
rect 161846 78920 161902 78976
rect 162214 79464 162270 79520
rect 162214 78784 162270 78840
rect 162858 79736 162914 79792
rect 162490 79600 162546 79656
rect 162306 76472 162362 76528
rect 162766 79600 162822 79656
rect 162674 79464 162730 79520
rect 162582 75928 162638 75984
rect 163226 79636 163228 79656
rect 163228 79636 163280 79656
rect 163280 79636 163282 79656
rect 163916 79872 163972 79928
rect 164376 79872 164432 79928
rect 163226 79600 163282 79636
rect 163502 79192 163558 79248
rect 163318 76064 163374 76120
rect 163778 79620 163834 79656
rect 164422 79736 164478 79792
rect 164744 79872 164800 79928
rect 163778 79600 163780 79620
rect 163780 79600 163832 79620
rect 163832 79600 163834 79620
rect 164238 79620 164294 79656
rect 163686 75928 163742 75984
rect 164238 79600 164240 79620
rect 164240 79600 164292 79620
rect 164292 79600 164294 79620
rect 164054 79464 164110 79520
rect 164054 71440 164110 71496
rect 164698 79736 164754 79792
rect 164928 79756 164984 79792
rect 164928 79736 164930 79756
rect 164930 79736 164982 79756
rect 164982 79736 164984 79756
rect 165296 79872 165352 79928
rect 164790 79464 164846 79520
rect 165066 77560 165122 77616
rect 164974 76064 165030 76120
rect 165664 79906 165720 79962
rect 166032 79872 166088 79928
rect 166584 79872 166640 79928
rect 165250 79192 165306 79248
rect 165894 79736 165950 79792
rect 165526 79600 165582 79656
rect 161294 4800 161350 4856
rect 165710 79056 165766 79112
rect 166446 75928 166502 75984
rect 166952 79872 167008 79928
rect 167136 79872 167192 79928
rect 167320 79838 167376 79894
rect 167504 79872 167560 79928
rect 166630 79636 166632 79656
rect 166632 79636 166684 79656
rect 166684 79636 166686 79656
rect 166630 79600 166686 79636
rect 166630 78512 166686 78568
rect 166722 77968 166778 78024
rect 166814 75928 166870 75984
rect 167090 79600 167146 79656
rect 166998 79192 167054 79248
rect 167274 79600 167330 79656
rect 167780 79906 167836 79962
rect 167550 79600 167606 79656
rect 167458 79464 167514 79520
rect 167366 79056 167422 79112
rect 167550 79056 167606 79112
rect 168056 79872 168112 79928
rect 168240 79906 168296 79962
rect 168424 79824 168480 79826
rect 168424 79772 168426 79824
rect 168426 79772 168478 79824
rect 168478 79772 168480 79824
rect 168424 79770 168480 79772
rect 168010 79600 168066 79656
rect 168010 79500 168012 79520
rect 168012 79500 168064 79520
rect 168064 79500 168066 79520
rect 168010 79464 168066 79500
rect 168792 79872 168848 79928
rect 169160 79906 169216 79962
rect 168378 79464 168434 79520
rect 168286 78648 168342 78704
rect 168194 75928 168250 75984
rect 169022 79736 169078 79792
rect 168562 77696 168618 77752
rect 169022 79192 169078 79248
rect 168930 78240 168986 78296
rect 169436 79906 169492 79962
rect 170080 79906 170136 79962
rect 169206 79464 169262 79520
rect 169390 79620 169446 79656
rect 169390 79600 169392 79620
rect 169392 79600 169444 79620
rect 169444 79600 169446 79620
rect 170448 79872 170504 79928
rect 169390 79328 169446 79384
rect 169114 76880 169170 76936
rect 169758 79056 169814 79112
rect 170310 79328 170366 79384
rect 170218 76472 170274 76528
rect 170494 79056 170550 79112
rect 170494 78920 170550 78976
rect 171276 79872 171332 79928
rect 171000 79736 171056 79792
rect 171552 79872 171608 79928
rect 170862 79636 170864 79656
rect 170864 79636 170916 79656
rect 170916 79636 170918 79656
rect 170862 79600 170918 79636
rect 170770 77560 170826 77616
rect 170770 76608 170826 76664
rect 171046 79464 171102 79520
rect 171230 78920 171286 78976
rect 171322 77968 171378 78024
rect 171506 79192 171562 79248
rect 172104 79872 172160 79928
rect 171874 79600 171930 79656
rect 171690 79464 171746 79520
rect 171690 79192 171746 79248
rect 171874 78240 171930 78296
rect 171598 76472 171654 76528
rect 171782 26968 171838 27024
rect 172288 79872 172344 79928
rect 172058 79464 172114 79520
rect 171966 77832 172022 77888
rect 172748 79906 172804 79962
rect 172932 79960 172988 79962
rect 172932 79908 172934 79960
rect 172934 79908 172986 79960
rect 172986 79908 172988 79960
rect 172932 79906 172988 79908
rect 172334 79192 172390 79248
rect 172242 78920 172298 78976
rect 172058 77560 172114 77616
rect 172426 78512 172482 78568
rect 173484 79872 173540 79928
rect 173852 79906 173908 79962
rect 173254 79600 173310 79656
rect 173254 79464 173310 79520
rect 173070 79192 173126 79248
rect 173346 79056 173402 79112
rect 173714 79464 173770 79520
rect 173714 78512 173770 78568
rect 173806 75928 173862 75984
rect 174312 79872 174368 79928
rect 174082 79464 174138 79520
rect 174542 79736 174598 79792
rect 175232 79872 175288 79928
rect 174082 75656 174138 75712
rect 173898 74296 173954 74352
rect 174542 75384 174598 75440
rect 175140 79736 175196 79792
rect 175416 79872 175472 79928
rect 175784 79872 175840 79928
rect 174818 79636 174820 79656
rect 174820 79636 174872 79656
rect 174872 79636 174874 79656
rect 174818 79600 174874 79636
rect 174818 78512 174874 78568
rect 174726 75520 174782 75576
rect 174726 75384 174782 75440
rect 175278 79620 175334 79656
rect 175278 79600 175280 79620
rect 175280 79600 175332 79620
rect 175332 79600 175334 79620
rect 175186 79464 175242 79520
rect 175186 78240 175242 78296
rect 175094 77016 175150 77072
rect 175002 76880 175058 76936
rect 174910 74296 174966 74352
rect 175186 73888 175242 73944
rect 176336 79872 176392 79928
rect 176198 79756 176254 79792
rect 176198 79736 176200 79756
rect 176200 79736 176252 79756
rect 176252 79736 176254 79756
rect 175462 73888 175518 73944
rect 175738 78920 175794 78976
rect 175646 72800 175702 72856
rect 175922 79464 175978 79520
rect 176520 79736 176576 79792
rect 176106 79620 176162 79656
rect 176106 79600 176108 79620
rect 176108 79600 176160 79620
rect 176160 79600 176162 79620
rect 176014 78104 176070 78160
rect 176290 77152 176346 77208
rect 176658 79464 176714 79520
rect 176566 75520 176622 75576
rect 176474 72800 176530 72856
rect 176842 78240 176898 78296
rect 177348 79906 177404 79962
rect 177532 79906 177588 79962
rect 177486 79736 177542 79792
rect 177210 77868 177212 77888
rect 177212 77868 177264 77888
rect 177264 77868 177266 77888
rect 177210 77832 177266 77868
rect 177670 79464 177726 79520
rect 177578 79192 177634 79248
rect 177854 78240 177910 78296
rect 178038 77560 178094 77616
rect 181442 80416 181498 80472
rect 181442 80144 181498 80200
rect 179326 80008 179382 80064
rect 178590 76880 178646 76936
rect 178038 72392 178094 72448
rect 179234 77832 179290 77888
rect 181074 79464 181130 79520
rect 179510 78920 179566 78976
rect 180890 78920 180946 78976
rect 182086 79736 182142 79792
rect 181166 78920 181222 78976
rect 179326 77152 179382 77208
rect 180062 77152 180118 77208
rect 181534 77868 181536 77888
rect 181536 77868 181588 77888
rect 181588 77868 181590 77888
rect 181534 77832 181590 77868
rect 182086 77424 182142 77480
rect 182914 69944 182970 70000
rect 183006 68856 183062 68912
rect 183558 74976 183614 75032
rect 185582 77424 185638 77480
rect 184202 68312 184258 68368
rect 186870 80144 186926 80200
rect 186686 76472 186742 76528
rect 187330 139168 187386 139224
rect 187514 138216 187570 138272
rect 187422 138080 187478 138136
rect 187422 80144 187478 80200
rect 187330 75792 187386 75848
rect 187698 77424 187754 77480
rect 187422 69672 187478 69728
rect 186962 62056 187018 62112
rect 186594 57840 186650 57896
rect 189078 200640 189134 200696
rect 188250 139304 188306 139360
rect 188066 75112 188122 75168
rect 187882 66136 187938 66192
rect 187882 65864 187938 65920
rect 187790 63144 187846 63200
rect 188526 127608 188582 127664
rect 188434 80416 188490 80472
rect 188434 71304 188490 71360
rect 189446 259528 189502 259584
rect 189538 143248 189594 143304
rect 189814 139712 189870 139768
rect 189170 67496 189226 67552
rect 189722 68176 189778 68232
rect 189354 67360 189410 67416
rect 189078 63008 189134 63064
rect 188250 59064 188306 59120
rect 189906 67360 189962 67416
rect 189906 66952 189962 67008
rect 191010 262248 191066 262304
rect 191838 262248 191894 262304
rect 190918 142976 190974 143032
rect 191378 259936 191434 259992
rect 190826 140700 190828 140720
rect 190828 140700 190880 140720
rect 190880 140700 190882 140720
rect 190826 140664 190882 140700
rect 190826 138624 190882 138680
rect 190642 61920 190698 61976
rect 190550 57568 190606 57624
rect 191102 138488 191158 138544
rect 191378 143112 191434 143168
rect 191470 74432 191526 74488
rect 191470 73752 191526 73808
rect 191746 61920 191802 61976
rect 191746 61512 191802 61568
rect 190826 56344 190882 56400
rect 192298 138352 192354 138408
rect 193402 144880 193458 144936
rect 193402 138896 193458 138952
rect 191930 58792 191986 58848
rect 191838 54984 191894 55040
rect 191838 54712 191894 54768
rect 190458 50768 190514 50824
rect 193586 66000 193642 66056
rect 193862 66816 193918 66872
rect 193770 57432 193826 57488
rect 193402 54848 193458 54904
rect 193402 54576 193458 54632
rect 194506 66000 194562 66056
rect 194506 65728 194562 65784
rect 194966 139032 195022 139088
rect 195334 146920 195390 146976
rect 195334 81232 195390 81288
rect 195058 79056 195114 79112
rect 195518 81096 195574 81152
rect 194782 53624 194838 53680
rect 194782 53216 194838 53272
rect 194690 52264 194746 52320
rect 194690 51856 194746 51912
rect 196530 137944 196586 138000
rect 197082 80960 197138 81016
rect 196162 66680 196218 66736
rect 196070 62056 196126 62112
rect 196162 58656 196218 58712
rect 195978 49408 196034 49464
rect 195978 49000 196034 49056
rect 194598 47640 194654 47696
rect 194598 44920 194654 44976
rect 197358 56208 197414 56264
rect 234618 278024 234674 278080
rect 299478 276664 299534 276720
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580262 365064 580318 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 477498 262792 477554 262848
rect 198738 196832 198794 196888
rect 198094 146240 198150 146296
rect 198094 137808 198150 137864
rect 198002 78920 198058 78976
rect 197450 55120 197506 55176
rect 197450 54440 197506 54496
rect 200302 200232 200358 200288
rect 200118 196696 200174 196752
rect 199106 80824 199162 80880
rect 199382 68876 199438 68912
rect 199382 68856 199384 68876
rect 199384 68856 199436 68876
rect 199436 68856 199438 68876
rect 199014 61784 199070 61840
rect 199014 61376 199070 61432
rect 198922 60560 198978 60616
rect 198830 57296 198886 57352
rect 198738 50904 198794 50960
rect 199566 50904 199622 50960
rect 199566 50224 199622 50280
rect 200210 196560 200266 196616
rect 201774 200096 201830 200152
rect 200302 63416 200358 63472
rect 200210 53760 200266 53816
rect 200118 49544 200174 49600
rect 201038 147736 201094 147792
rect 200762 69536 200818 69592
rect 200670 44104 200726 44160
rect 201406 63416 201462 63472
rect 201406 62872 201462 62928
rect 201406 53760 201462 53816
rect 201406 53080 201462 53136
rect 201406 49544 201462 49600
rect 201406 48864 201462 48920
rect 201682 55156 201684 55176
rect 201684 55156 201736 55176
rect 201736 55156 201738 55176
rect 201682 55120 201738 55156
rect 201866 59200 201922 59256
rect 202786 59200 202842 59256
rect 202786 58520 202842 58576
rect 201958 56480 202014 56536
rect 202786 56480 202842 56536
rect 202786 56072 202842 56128
rect 201774 52400 201830 52456
rect 202786 52400 202842 52456
rect 202786 51720 202842 51776
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580446 232328 580502 232384
rect 580354 219000 580410 219056
rect 579802 205672 579858 205728
rect 205730 193024 205786 193080
rect 204258 192616 204314 192672
rect 203154 77288 203210 77344
rect 203062 50904 203118 50960
rect 203706 78240 203762 78296
rect 203614 68176 203670 68232
rect 203338 48184 203394 48240
rect 202878 43968 202934 44024
rect 202878 43424 202934 43480
rect 204166 77968 204222 78024
rect 204166 77288 204222 77344
rect 204258 55936 204314 55992
rect 204166 48184 204222 48240
rect 204166 47504 204222 47560
rect 204626 76608 204682 76664
rect 205914 192888 205970 192944
rect 205822 192480 205878 192536
rect 206006 192752 206062 192808
rect 205914 76880 205970 76936
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580354 152632 580410 152688
rect 289082 139576 289138 139632
rect 205914 76472 205970 76528
rect 211802 76744 211858 76800
rect 206190 75656 206246 75712
rect 206558 75656 206614 75712
rect 206558 75112 206614 75168
rect 205638 73072 205694 73128
rect 205638 72392 205694 72448
rect 213918 67088 213974 67144
rect 212538 32408 212594 32464
rect 227718 63280 227774 63336
rect 231858 61648 231914 61704
rect 230478 42064 230534 42120
rect 229098 18536 229154 18592
rect 247682 76608 247738 76664
rect 242898 67224 242954 67280
rect 249798 44784 249854 44840
rect 269762 77968 269818 78024
rect 263598 57704 263654 57760
rect 267738 40568 267794 40624
rect 264978 26832 265034 26888
rect 287702 77832 287758 77888
rect 274638 65864 274694 65920
rect 277398 63144 277454 63200
rect 281538 58928 281594 58984
rect 284390 53352 284446 53408
rect 295338 66952 295394 67008
rect 292578 63008 292634 63064
rect 304998 73752 305054 73808
rect 301502 72392 301558 72448
rect 309138 61512 309194 61568
rect 313278 57568 313334 57624
rect 576122 139440 576178 139496
rect 523130 80824 523186 80880
rect 327078 58792 327134 58848
rect 331218 54712 331274 54768
rect 338118 50360 338174 50416
rect 336278 11600 336334 11656
rect 349158 56344 349214 56400
rect 356058 49136 356114 49192
rect 382278 78784 382334 78840
rect 362958 65728 363014 65784
rect 364982 57432 365038 57488
rect 376758 66816 376814 66872
rect 369858 54576 369914 54632
rect 373998 47640 374054 47696
rect 380898 58656 380954 58712
rect 436098 78648 436154 78704
rect 382922 53216 382978 53272
rect 387798 49000 387854 49056
rect 398838 56208 398894 56264
rect 412638 60016 412694 60072
rect 401598 54440 401654 54496
rect 405738 51856 405794 51912
rect 414662 57296 414718 57352
rect 418802 50224 418858 50280
rect 422942 61376 422998 61432
rect 427818 43560 427874 43616
rect 430578 62872 430634 62928
rect 453302 75248 453358 75304
rect 437478 53080 437534 53136
rect 440238 48864 440294 48920
rect 450542 58520 450598 58576
rect 459558 56072 459614 56128
rect 455418 51720 455474 51776
rect 458178 46144 458234 46200
rect 470598 47504 470654 47560
rect 476118 43424 476174 43480
rect 489182 71304 489238 71360
rect 498198 69672 498254 69728
rect 494058 36488 494114 36544
rect 499578 55936 499634 55992
rect 507858 71168 507914 71224
rect 514022 65592 514078 65648
rect 511998 64232 512054 64288
rect 525798 80688 525854 80744
rect 536838 78920 536894 78976
rect 535458 75112 535514 75168
rect 531318 71032 531374 71088
rect 527822 65456 527878 65512
rect 553398 76472 553454 76528
rect 543738 64096 543794 64152
rect 547878 62736 547934 62792
rect 545762 57160 545818 57216
rect 561678 69536 561734 69592
rect 565818 68176 565874 68232
rect 563702 55800 563758 55856
rect 567842 59880 567898 59936
rect 580446 139304 580502 139360
rect 580262 99456 580318 99512
rect 580170 86128 580226 86184
rect 580998 78512 581054 78568
rect 580170 72936 580226 72992
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2773 371378 2839 371381
rect -960 371376 2839 371378
rect -960 371320 2778 371376
rect 2834 371320 2839 371376
rect -960 371318 2839 371320
rect -960 371228 480 371318
rect 2773 371315 2839 371318
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 189022 278020 189028 278084
rect 189092 278082 189098 278084
rect 234613 278082 234679 278085
rect 189092 278080 234679 278082
rect 189092 278024 234618 278080
rect 234674 278024 234679 278080
rect 189092 278022 234679 278024
rect 189092 278020 189098 278022
rect 234613 278019 234679 278022
rect 156045 277538 156111 277541
rect 189022 277538 189028 277540
rect 156045 277536 189028 277538
rect 156045 277480 156050 277536
rect 156106 277480 189028 277536
rect 156045 277478 189028 277480
rect 156045 277475 156111 277478
rect 189022 277476 189028 277478
rect 189092 277476 189098 277540
rect 299473 276722 299539 276725
rect 190410 276720 299539 276722
rect 190410 276664 299478 276720
rect 299534 276664 299539 276720
rect 190410 276662 299539 276664
rect 153377 276042 153443 276045
rect 189206 276042 189212 276044
rect 153377 276040 189212 276042
rect 153377 275984 153382 276040
rect 153438 275984 189212 276040
rect 153377 275982 189212 275984
rect 153377 275979 153443 275982
rect 189206 275980 189212 275982
rect 189276 276042 189282 276044
rect 190410 276042 190470 276662
rect 299473 276659 299539 276662
rect 189276 275982 190470 276042
rect 189276 275980 189282 275982
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 162209 265570 162275 265573
rect 167453 265570 167519 265573
rect 162209 265568 167519 265570
rect 162209 265512 162214 265568
rect 162270 265512 167458 265568
rect 167514 265512 167519 265568
rect 162209 265510 167519 265512
rect 162209 265507 162275 265510
rect 167453 265507 167519 265510
rect 167545 265434 167611 265437
rect 197486 265434 197492 265436
rect 167545 265432 197492 265434
rect 167545 265376 167550 265432
rect 167606 265376 197492 265432
rect 167545 265374 197492 265376
rect 167545 265371 167611 265374
rect 197486 265372 197492 265374
rect 197556 265372 197562 265436
rect 165153 265298 165219 265301
rect 196198 265298 196204 265300
rect 165153 265296 196204 265298
rect 165153 265240 165158 265296
rect 165214 265240 196204 265296
rect 165153 265238 196204 265240
rect 165153 265235 165219 265238
rect 196198 265236 196204 265238
rect 196268 265236 196274 265300
rect 111558 265100 111564 265164
rect 111628 265162 111634 265164
rect 135897 265162 135963 265165
rect 111628 265160 135963 265162
rect 111628 265104 135902 265160
rect 135958 265104 135963 265160
rect 111628 265102 135963 265104
rect 111628 265100 111634 265102
rect 135897 265099 135963 265102
rect 163497 265162 163563 265165
rect 167453 265162 167519 265165
rect 194542 265162 194548 265164
rect 163497 265160 167378 265162
rect 163497 265104 163502 265160
rect 163558 265104 167378 265160
rect 163497 265102 167378 265104
rect 163497 265099 163563 265102
rect 113030 264964 113036 265028
rect 113100 265026 113106 265028
rect 138749 265026 138815 265029
rect 113100 265024 138815 265026
rect 113100 264968 138754 265024
rect 138810 264968 138815 265024
rect 113100 264966 138815 264968
rect 113100 264964 113106 264966
rect 138749 264963 138815 264966
rect 164877 265026 164943 265029
rect 165153 265026 165219 265029
rect 164877 265024 165219 265026
rect 164877 264968 164882 265024
rect 164938 264968 165158 265024
rect 165214 264968 165219 265024
rect 164877 264966 165219 264968
rect 167318 265026 167378 265102
rect 167453 265160 194548 265162
rect 167453 265104 167458 265160
rect 167514 265104 194548 265160
rect 167453 265102 194548 265104
rect 167453 265099 167519 265102
rect 194542 265100 194548 265102
rect 194612 265100 194618 265164
rect 197670 265026 197676 265028
rect 167318 264966 197676 265026
rect 164877 264963 164943 264966
rect 165153 264963 165219 264966
rect 197670 264964 197676 264966
rect 197740 264964 197746 265028
rect 119838 263876 119844 263940
rect 119908 263938 119914 263940
rect 146201 263938 146267 263941
rect 119908 263936 146267 263938
rect 119908 263880 146206 263936
rect 146262 263880 146267 263936
rect 119908 263878 146267 263880
rect 119908 263876 119914 263878
rect 146201 263875 146267 263878
rect 121310 263740 121316 263804
rect 121380 263802 121386 263804
rect 147765 263802 147831 263805
rect 121380 263800 147831 263802
rect 121380 263744 147770 263800
rect 147826 263744 147831 263800
rect 121380 263742 147831 263744
rect 121380 263740 121386 263742
rect 147765 263739 147831 263742
rect 112846 263604 112852 263668
rect 112916 263666 112922 263668
rect 145281 263666 145347 263669
rect 145557 263666 145623 263669
rect 112916 263664 145623 263666
rect 112916 263608 145286 263664
rect 145342 263608 145562 263664
rect 145618 263608 145623 263664
rect 112916 263606 145623 263608
rect 112916 263604 112922 263606
rect 145281 263603 145347 263606
rect 145557 263603 145623 263606
rect 163405 263258 163471 263261
rect 163589 263258 163655 263261
rect 163405 263256 163655 263258
rect 163405 263200 163410 263256
rect 163466 263200 163594 263256
rect 163650 263200 163655 263256
rect 163405 263198 163655 263200
rect 163405 263195 163471 263198
rect 163589 263195 163655 263198
rect 114134 262924 114140 262988
rect 114204 262986 114210 262988
rect 148501 262986 148567 262989
rect 114204 262984 148567 262986
rect 114204 262928 148506 262984
rect 148562 262928 148567 262984
rect 114204 262926 148567 262928
rect 114204 262924 114210 262926
rect 148501 262923 148567 262926
rect 115606 262788 115612 262852
rect 115676 262850 115682 262852
rect 138657 262850 138723 262853
rect 477493 262850 477559 262853
rect 115676 262848 138723 262850
rect 115676 262792 138662 262848
rect 138718 262792 138723 262848
rect 115676 262790 138723 262792
rect 115676 262788 115682 262790
rect 138657 262787 138723 262790
rect 151770 262848 477559 262850
rect 151770 262792 477498 262848
rect 477554 262792 477559 262848
rect 151770 262790 477559 262792
rect 112662 262652 112668 262716
rect 112732 262714 112738 262716
rect 140313 262714 140379 262717
rect 112732 262712 140379 262714
rect 112732 262656 140318 262712
rect 140374 262656 140379 262712
rect 112732 262654 140379 262656
rect 112732 262652 112738 262654
rect 140313 262651 140379 262654
rect 113950 262516 113956 262580
rect 114020 262578 114026 262580
rect 146937 262578 147003 262581
rect 114020 262576 147003 262578
rect 114020 262520 146942 262576
rect 146998 262520 147003 262576
rect 114020 262518 147003 262520
rect 114020 262516 114026 262518
rect 146937 262515 147003 262518
rect 116710 262380 116716 262444
rect 116780 262442 116786 262444
rect 150525 262442 150591 262445
rect 151770 262442 151830 262790
rect 477493 262787 477559 262790
rect 158805 262714 158871 262717
rect 159909 262714 159975 262717
rect 193438 262714 193444 262716
rect 158805 262712 193444 262714
rect 158805 262656 158810 262712
rect 158866 262656 159914 262712
rect 159970 262656 193444 262712
rect 158805 262654 193444 262656
rect 158805 262651 158871 262654
rect 159909 262651 159975 262654
rect 193438 262652 193444 262654
rect 193508 262652 193514 262716
rect 163405 262578 163471 262581
rect 191966 262578 191972 262580
rect 163405 262576 191972 262578
rect 163405 262520 163410 262576
rect 163466 262520 191972 262576
rect 163405 262518 191972 262520
rect 163405 262515 163471 262518
rect 191966 262516 191972 262518
rect 192036 262516 192042 262580
rect 116780 262440 151830 262442
rect 116780 262384 150530 262440
rect 150586 262384 151830 262440
rect 116780 262382 151830 262384
rect 162025 262442 162091 262445
rect 193622 262442 193628 262444
rect 162025 262440 193628 262442
rect 162025 262384 162030 262440
rect 162086 262384 193628 262440
rect 162025 262382 193628 262384
rect 116780 262380 116786 262382
rect 150525 262379 150591 262382
rect 162025 262379 162091 262382
rect 193622 262380 193628 262382
rect 193692 262380 193698 262444
rect 115422 262244 115428 262308
rect 115492 262306 115498 262308
rect 129825 262306 129891 262309
rect 115492 262304 129891 262306
rect 115492 262248 129830 262304
rect 129886 262248 129891 262304
rect 115492 262246 129891 262248
rect 115492 262244 115498 262246
rect 129825 262243 129891 262246
rect 190494 262244 190500 262308
rect 190564 262306 190570 262308
rect 191005 262306 191071 262309
rect 190564 262304 191071 262306
rect 190564 262248 191010 262304
rect 191066 262248 191071 262304
rect 190564 262246 191071 262248
rect 190564 262244 190570 262246
rect 191005 262243 191071 262246
rect 191833 262306 191899 262309
rect 192150 262306 192156 262308
rect 191833 262304 192156 262306
rect 191833 262248 191838 262304
rect 191894 262248 192156 262304
rect 191833 262246 192156 262248
rect 191833 262243 191899 262246
rect 192150 262244 192156 262246
rect 192220 262244 192226 262308
rect 111374 261020 111380 261084
rect 111444 261082 111450 261084
rect 132033 261082 132099 261085
rect 111444 261080 132099 261082
rect 111444 261024 132038 261080
rect 132094 261024 132099 261080
rect 111444 261022 132099 261024
rect 111444 261020 111450 261022
rect 132033 261019 132099 261022
rect 111190 260884 111196 260948
rect 111260 260946 111266 260948
rect 137461 260946 137527 260949
rect 111260 260944 137527 260946
rect 111260 260888 137466 260944
rect 137522 260888 137527 260944
rect 111260 260886 137527 260888
rect 111260 260884 111266 260886
rect 137461 260883 137527 260886
rect 161473 260810 161539 260813
rect 162669 260810 162735 260813
rect 161473 260808 162735 260810
rect 161473 260752 161478 260808
rect 161534 260752 162674 260808
rect 162730 260752 162735 260808
rect 161473 260750 162735 260752
rect 161473 260747 161539 260750
rect 162669 260747 162735 260750
rect 117078 260340 117084 260404
rect 117148 260402 117154 260404
rect 139669 260402 139735 260405
rect 117148 260400 139735 260402
rect 117148 260344 139674 260400
rect 139730 260344 139735 260400
rect 117148 260342 139735 260344
rect 117148 260340 117154 260342
rect 139669 260339 139735 260342
rect 121126 260204 121132 260268
rect 121196 260266 121202 260268
rect 143625 260266 143691 260269
rect 144499 260266 144565 260269
rect 121196 260264 144565 260266
rect 121196 260208 143630 260264
rect 143686 260208 144504 260264
rect 144560 260208 144565 260264
rect 121196 260206 144565 260208
rect 121196 260204 121202 260206
rect 143625 260203 143691 260206
rect 144499 260203 144565 260206
rect 157333 260266 157399 260269
rect 158299 260266 158365 260269
rect 157333 260264 158365 260266
rect 157333 260208 157338 260264
rect 157394 260208 158304 260264
rect 158360 260208 158365 260264
rect 157333 260206 158365 260208
rect 157333 260203 157399 260206
rect 158299 260203 158365 260206
rect 118366 260068 118372 260132
rect 118436 260130 118442 260132
rect 140773 260130 140839 260133
rect 141739 260130 141805 260133
rect 142429 260130 142495 260133
rect 143395 260130 143461 260133
rect 189574 260130 189580 260132
rect 118436 260128 141805 260130
rect 118436 260072 140778 260128
rect 140834 260072 141744 260128
rect 141800 260072 141805 260128
rect 118436 260070 141805 260072
rect 118436 260068 118442 260070
rect 140773 260067 140839 260070
rect 141739 260067 141805 260070
rect 142110 260128 143461 260130
rect 142110 260072 142434 260128
rect 142490 260072 143400 260128
rect 143456 260072 143461 260128
rect 142110 260070 143461 260072
rect 116894 259932 116900 259996
rect 116964 259994 116970 259996
rect 142110 259994 142170 260070
rect 142429 260067 142495 260070
rect 143395 260067 143461 260070
rect 180750 260070 189580 260130
rect 116964 259934 142170 259994
rect 160093 259994 160159 259997
rect 160921 259994 160987 259997
rect 180750 259994 180810 260070
rect 189574 260068 189580 260070
rect 189644 260068 189650 260132
rect 191373 259994 191439 259997
rect 160093 259992 180810 259994
rect 160093 259936 160098 259992
rect 160154 259936 160926 259992
rect 160982 259936 180810 259992
rect 160093 259934 180810 259936
rect 185534 259992 191439 259994
rect 185534 259936 191378 259992
rect 191434 259936 191439 259992
rect 185534 259934 191439 259936
rect 116964 259932 116970 259934
rect 160093 259931 160159 259934
rect 160921 259931 160987 259934
rect 118182 259796 118188 259860
rect 118252 259858 118258 259860
rect 144913 259858 144979 259861
rect 118252 259856 144979 259858
rect 118252 259800 144918 259856
rect 144974 259800 144979 259856
rect 118252 259798 144979 259800
rect 118252 259796 118258 259798
rect 144913 259795 144979 259798
rect 162577 259858 162643 259861
rect 185534 259858 185594 259934
rect 191373 259931 191439 259934
rect 162577 259856 185594 259858
rect 162577 259800 162582 259856
rect 162638 259800 185594 259856
rect 162577 259798 185594 259800
rect 162577 259795 162643 259798
rect 113766 259660 113772 259724
rect 113836 259722 113842 259724
rect 146477 259722 146543 259725
rect 113836 259720 146543 259722
rect 113836 259664 146482 259720
rect 146538 259664 146543 259720
rect 113836 259662 146543 259664
rect 113836 259660 113842 259662
rect 146477 259659 146543 259662
rect 158621 259722 158687 259725
rect 191782 259722 191788 259724
rect 158621 259720 191788 259722
rect 158621 259664 158626 259720
rect 158682 259664 191788 259720
rect 158621 259662 191788 259664
rect 158621 259659 158687 259662
rect 191782 259660 191788 259662
rect 191852 259660 191858 259724
rect 115790 259524 115796 259588
rect 115860 259586 115866 259588
rect 149053 259586 149119 259589
rect 149789 259586 149855 259589
rect 115860 259584 149855 259586
rect 115860 259528 149058 259584
rect 149114 259528 149794 259584
rect 149850 259528 149855 259584
rect 115860 259526 149855 259528
rect 115860 259524 115866 259526
rect 149053 259523 149119 259526
rect 149789 259523 149855 259526
rect 155217 259586 155283 259589
rect 185669 259586 185735 259589
rect 186078 259586 186084 259588
rect 155217 259584 185594 259586
rect 155217 259528 155222 259584
rect 155278 259528 185594 259584
rect 155217 259526 185594 259528
rect 155217 259523 155283 259526
rect 185534 259450 185594 259526
rect 185669 259584 186084 259586
rect 185669 259528 185674 259584
rect 185730 259528 186084 259584
rect 185669 259526 186084 259528
rect 185669 259523 185735 259526
rect 186078 259524 186084 259526
rect 186148 259524 186154 259588
rect 189441 259586 189507 259589
rect 186270 259584 189507 259586
rect 186270 259528 189446 259584
rect 189502 259528 189507 259584
rect 186270 259526 189507 259528
rect 186270 259450 186330 259526
rect 189441 259523 189507 259526
rect 185534 259390 186330 259450
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 580441 232386 580507 232389
rect 583520 232386 584960 232476
rect 580441 232384 584960 232386
rect 580441 232328 580446 232384
rect 580502 232328 584960 232384
rect 580441 232326 584960 232328
rect 580441 232323 580507 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 186078 212468 186084 212532
rect 186148 212530 186154 212532
rect 187182 212530 187188 212532
rect 186148 212470 187188 212530
rect 186148 212468 186154 212470
rect 187182 212468 187188 212470
rect 187252 212468 187258 212532
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 119981 200698 120047 200701
rect 132033 200698 132099 200701
rect 119981 200696 132099 200698
rect 119981 200640 119986 200696
rect 120042 200640 132038 200696
rect 132094 200640 132099 200696
rect 119981 200638 132099 200640
rect 119981 200635 120047 200638
rect 132033 200635 132099 200638
rect 132217 200698 132283 200701
rect 141550 200698 141556 200700
rect 132217 200696 141556 200698
rect 132217 200640 132222 200696
rect 132278 200640 141556 200696
rect 132217 200638 141556 200640
rect 132217 200635 132283 200638
rect 141550 200636 141556 200638
rect 141620 200636 141626 200700
rect 178677 200698 178743 200701
rect 189073 200698 189139 200701
rect 178677 200696 189139 200698
rect 178677 200640 178682 200696
rect 178738 200640 189078 200696
rect 189134 200640 189139 200696
rect 178677 200638 189139 200640
rect 178677 200635 178743 200638
rect 189073 200635 189139 200638
rect 107377 200562 107443 200565
rect 136582 200562 136588 200564
rect 107377 200560 136588 200562
rect 107377 200504 107382 200560
rect 107438 200504 136588 200560
rect 107377 200502 136588 200504
rect 107377 200499 107443 200502
rect 136582 200500 136588 200502
rect 136652 200500 136658 200564
rect 107285 200426 107351 200429
rect 130469 200426 130535 200429
rect 107285 200424 130535 200426
rect 107285 200368 107290 200424
rect 107346 200368 130474 200424
rect 130530 200368 130535 200424
rect 107285 200366 130535 200368
rect 107285 200363 107351 200366
rect 130469 200363 130535 200366
rect 131297 200426 131363 200429
rect 138054 200426 138060 200428
rect 131297 200424 138060 200426
rect 131297 200368 131302 200424
rect 131358 200368 138060 200424
rect 131297 200366 138060 200368
rect 131297 200363 131363 200366
rect 138054 200364 138060 200366
rect 138124 200364 138130 200428
rect 127617 200290 127683 200293
rect 150198 200290 150204 200292
rect 127617 200288 150204 200290
rect 127617 200232 127622 200288
rect 127678 200232 150204 200288
rect 127617 200230 150204 200232
rect 127617 200227 127683 200230
rect 150198 200228 150204 200230
rect 150268 200228 150274 200292
rect 170254 200228 170260 200292
rect 170324 200290 170330 200292
rect 200297 200290 200363 200293
rect 170324 200288 200363 200290
rect 170324 200232 200302 200288
rect 200358 200232 200363 200288
rect 170324 200230 200363 200232
rect 170324 200228 170330 200230
rect 200297 200227 200363 200230
rect 130009 200154 130075 200157
rect 131297 200154 131363 200157
rect 130009 200152 131363 200154
rect 130009 200096 130014 200152
rect 130070 200096 131302 200152
rect 131358 200096 131363 200152
rect 130009 200094 131363 200096
rect 130009 200091 130075 200094
rect 131297 200091 131363 200094
rect 131665 200154 131731 200157
rect 133638 200154 133644 200156
rect 131665 200152 133644 200154
rect 131665 200096 131670 200152
rect 131726 200096 133644 200152
rect 131665 200094 133644 200096
rect 131665 200091 131731 200094
rect 133638 200092 133644 200094
rect 133708 200092 133714 200156
rect 138054 200092 138060 200156
rect 138124 200154 138130 200156
rect 138124 200094 142170 200154
rect 138124 200092 138130 200094
rect 132217 200018 132283 200021
rect 132217 200016 137754 200018
rect 132217 199960 132222 200016
rect 132278 199960 137754 200016
rect 132217 199958 137754 199960
rect 132217 199955 132283 199958
rect 137694 199885 137754 199958
rect 138606 199956 138612 200020
rect 138676 200018 138682 200020
rect 138676 199958 139226 200018
rect 138676 199956 138682 199958
rect 128997 199882 129063 199885
rect 131757 199882 131823 199885
rect 128997 199880 131823 199882
rect 128997 199824 129002 199880
rect 129058 199824 131762 199880
rect 131818 199824 131823 199880
rect 128997 199822 131823 199824
rect 128997 199819 129063 199822
rect 131757 199819 131823 199822
rect 132125 199882 132191 199885
rect 132907 199882 132973 199885
rect 132125 199880 132973 199882
rect 132125 199824 132130 199880
rect 132186 199824 132912 199880
rect 132968 199824 132973 199880
rect 132125 199822 132973 199824
rect 132125 199819 132191 199822
rect 132907 199819 132973 199822
rect 133086 199820 133092 199884
rect 133156 199882 133162 199884
rect 133367 199882 133433 199885
rect 133643 199884 133709 199885
rect 133638 199882 133644 199884
rect 133156 199880 133433 199882
rect 133156 199824 133372 199880
rect 133428 199824 133433 199880
rect 133156 199822 133433 199824
rect 133552 199822 133644 199882
rect 133156 199820 133162 199822
rect 133367 199819 133433 199822
rect 133638 199820 133644 199822
rect 133708 199820 133714 199884
rect 133919 199882 133985 199885
rect 134742 199882 134748 199884
rect 133919 199880 134748 199882
rect 133919 199824 133924 199880
rect 133980 199824 134748 199880
rect 133919 199822 134748 199824
rect 133643 199819 133709 199820
rect 133919 199819 133985 199822
rect 134742 199820 134748 199822
rect 134812 199820 134818 199884
rect 135483 199880 135549 199885
rect 135483 199824 135488 199880
rect 135544 199824 135549 199880
rect 135483 199819 135549 199824
rect 136030 199820 136036 199884
rect 136100 199882 136106 199884
rect 136495 199882 136561 199885
rect 136100 199880 136561 199882
rect 136100 199824 136500 199880
rect 136556 199824 136561 199880
rect 136100 199822 136561 199824
rect 136100 199820 136106 199822
rect 136495 199819 136561 199822
rect 136771 199880 136837 199885
rect 136771 199824 136776 199880
rect 136832 199824 136837 199880
rect 136771 199819 136837 199824
rect 137047 199882 137113 199885
rect 137047 199880 137386 199882
rect 137047 199824 137052 199880
rect 137108 199824 137386 199880
rect 137047 199822 137386 199824
rect 137047 199819 137113 199822
rect 135486 199749 135546 199819
rect 136774 199749 136834 199819
rect 131573 199746 131639 199749
rect 134425 199746 134491 199749
rect 131573 199744 134491 199746
rect 131573 199688 131578 199744
rect 131634 199688 134430 199744
rect 134486 199688 134491 199744
rect 131573 199686 134491 199688
rect 131573 199683 131639 199686
rect 134425 199683 134491 199686
rect 135437 199744 135546 199749
rect 135437 199688 135442 199744
rect 135498 199688 135546 199744
rect 135437 199686 135546 199688
rect 135437 199683 135503 199686
rect 136398 199684 136404 199748
rect 136468 199746 136474 199748
rect 136541 199746 136607 199749
rect 136468 199744 136607 199746
rect 136468 199688 136546 199744
rect 136602 199688 136607 199744
rect 136468 199686 136607 199688
rect 136774 199744 136883 199749
rect 136774 199688 136822 199744
rect 136878 199688 136883 199744
rect 136774 199686 136883 199688
rect 136468 199684 136474 199686
rect 136541 199683 136607 199686
rect 136817 199683 136883 199686
rect 137134 199684 137140 199748
rect 137204 199746 137210 199748
rect 137326 199746 137386 199822
rect 137691 199880 137757 199885
rect 137691 199824 137696 199880
rect 137752 199824 137757 199880
rect 137691 199819 137757 199824
rect 137875 199880 137941 199885
rect 137875 199824 137880 199880
rect 137936 199824 137941 199880
rect 137875 199819 137941 199824
rect 138059 199880 138125 199885
rect 138059 199824 138064 199880
rect 138120 199824 138125 199880
rect 138059 199819 138125 199824
rect 138243 199880 138309 199885
rect 138243 199824 138248 199880
rect 138304 199824 138309 199880
rect 138243 199819 138309 199824
rect 138427 199882 138493 199885
rect 138790 199882 138796 199884
rect 138427 199880 138796 199882
rect 138427 199824 138432 199880
rect 138488 199824 138796 199880
rect 138427 199822 138796 199824
rect 138427 199819 138493 199822
rect 138790 199820 138796 199822
rect 138860 199820 138866 199884
rect 138979 199882 139045 199885
rect 139166 199882 139226 199958
rect 142110 199919 142170 200094
rect 148182 200094 149576 200154
rect 148182 199919 148242 200094
rect 139439 199916 139505 199919
rect 138979 199880 139226 199882
rect 138979 199824 138984 199880
rect 139040 199824 139226 199880
rect 138979 199822 139226 199824
rect 139396 199914 139505 199916
rect 139396 199858 139444 199914
rect 139500 199858 139505 199914
rect 142107 199914 142173 199919
rect 139396 199853 139505 199858
rect 140083 199882 140149 199885
rect 141003 199884 141069 199885
rect 140630 199882 140636 199884
rect 140083 199880 140636 199882
rect 138979 199819 139045 199822
rect 137204 199686 137386 199746
rect 137204 199684 137210 199686
rect 137686 199684 137692 199748
rect 137756 199746 137762 199748
rect 137878 199746 137938 199819
rect 137756 199686 137938 199746
rect 137756 199684 137762 199686
rect 138062 199613 138122 199819
rect 138246 199613 138306 199819
rect 138933 199746 138999 199749
rect 139396 199746 139456 199853
rect 140083 199824 140088 199880
rect 140144 199824 140636 199880
rect 140083 199822 140636 199824
rect 140083 199819 140149 199822
rect 140630 199820 140636 199822
rect 140700 199820 140706 199884
rect 140998 199882 141004 199884
rect 140912 199822 141004 199882
rect 140998 199820 141004 199822
rect 141068 199820 141074 199884
rect 141279 199882 141345 199885
rect 141279 199880 141388 199882
rect 141279 199824 141284 199880
rect 141340 199824 141388 199880
rect 141003 199819 141069 199820
rect 141279 199819 141388 199824
rect 141555 199880 141621 199885
rect 141555 199824 141560 199880
rect 141616 199824 141621 199880
rect 142107 199858 142112 199914
rect 142168 199858 142173 199914
rect 142475 199914 142541 199919
rect 142475 199884 142480 199914
rect 142536 199884 142541 199914
rect 144499 199914 144565 199919
rect 142107 199853 142173 199858
rect 141555 199819 141621 199824
rect 142470 199820 142476 199884
rect 142540 199882 142546 199884
rect 142540 199822 142598 199882
rect 143487 199880 143553 199885
rect 144499 199884 144504 199914
rect 144560 199884 144565 199914
rect 145419 199914 145485 199919
rect 147535 199916 147601 199919
rect 145419 199884 145424 199914
rect 145480 199884 145485 199914
rect 147492 199914 147601 199916
rect 143487 199824 143492 199880
rect 143548 199824 143553 199880
rect 142540 199820 142546 199822
rect 143487 199819 143553 199824
rect 144494 199820 144500 199884
rect 144564 199882 144570 199884
rect 144564 199822 144622 199882
rect 144564 199820 144570 199822
rect 145414 199820 145420 199884
rect 145484 199882 145490 199884
rect 145484 199822 145542 199882
rect 146155 199880 146221 199885
rect 146155 199824 146160 199880
rect 146216 199824 146221 199880
rect 145484 199820 145490 199822
rect 146155 199819 146221 199824
rect 147070 199820 147076 199884
rect 147140 199882 147146 199884
rect 147492 199882 147540 199914
rect 147140 199858 147540 199882
rect 147596 199858 147601 199914
rect 147995 199914 148061 199919
rect 147811 199884 147877 199885
rect 147995 199884 148000 199914
rect 148056 199884 148061 199914
rect 148179 199914 148245 199919
rect 149375 199916 149441 199919
rect 147806 199882 147812 199884
rect 147140 199853 147601 199858
rect 147140 199822 147552 199853
rect 147720 199822 147812 199882
rect 147140 199820 147146 199822
rect 147806 199820 147812 199822
rect 147876 199820 147882 199884
rect 147990 199820 147996 199884
rect 148060 199882 148066 199884
rect 148060 199822 148118 199882
rect 148179 199858 148184 199914
rect 148240 199858 148245 199914
rect 149332 199914 149441 199916
rect 148179 199853 148245 199858
rect 148060 199820 148066 199822
rect 148542 199820 148548 199884
rect 148612 199882 148618 199884
rect 149332 199882 149380 199914
rect 148612 199858 149380 199882
rect 149436 199858 149441 199914
rect 148612 199853 149441 199858
rect 148612 199822 149392 199853
rect 148612 199820 148618 199822
rect 147811 199819 147877 199820
rect 140819 199748 140885 199749
rect 138933 199744 139456 199746
rect 138933 199688 138938 199744
rect 138994 199688 139456 199744
rect 138933 199686 139456 199688
rect 138933 199683 138999 199686
rect 140078 199684 140084 199748
rect 140148 199746 140154 199748
rect 140148 199715 140330 199746
rect 140148 199710 140333 199715
rect 140148 199686 140272 199710
rect 140148 199684 140154 199686
rect 140267 199654 140272 199686
rect 140328 199654 140333 199710
rect 140814 199684 140820 199748
rect 140884 199746 140890 199748
rect 140884 199686 140976 199746
rect 140884 199684 140890 199686
rect 140819 199683 140885 199684
rect 140267 199649 140333 199654
rect 141328 199613 141388 199819
rect 141558 199749 141618 199819
rect 141509 199744 141618 199749
rect 141509 199688 141514 199744
rect 141570 199688 141618 199744
rect 141509 199686 141618 199688
rect 143165 199746 143231 199749
rect 143490 199746 143550 199819
rect 143165 199744 143550 199746
rect 143165 199688 143170 199744
rect 143226 199688 143550 199744
rect 143165 199686 143550 199688
rect 141509 199683 141575 199686
rect 143165 199683 143231 199686
rect 145598 199684 145604 199748
rect 145668 199746 145674 199748
rect 146158 199746 146218 199819
rect 148409 199746 148475 199749
rect 145668 199686 146218 199746
rect 147814 199744 148475 199746
rect 147814 199688 148414 199744
rect 148470 199688 148475 199744
rect 147814 199686 148475 199688
rect 145668 199684 145674 199686
rect 106089 199610 106155 199613
rect 129549 199610 129615 199613
rect 106089 199608 129615 199610
rect 106089 199552 106094 199608
rect 106150 199552 129554 199608
rect 129610 199552 129615 199608
rect 106089 199550 129615 199552
rect 106089 199547 106155 199550
rect 129549 199547 129615 199550
rect 132493 199610 132559 199613
rect 136449 199610 136515 199613
rect 136633 199612 136699 199613
rect 132493 199608 136515 199610
rect 132493 199552 132498 199608
rect 132554 199552 136454 199608
rect 136510 199552 136515 199608
rect 132493 199550 136515 199552
rect 132493 199547 132559 199550
rect 136449 199547 136515 199550
rect 136582 199548 136588 199612
rect 136652 199610 136699 199612
rect 136652 199608 136744 199610
rect 136694 199552 136744 199608
rect 136652 199550 136744 199552
rect 138062 199608 138171 199613
rect 138062 199552 138110 199608
rect 138166 199552 138171 199608
rect 138062 199550 138171 199552
rect 138246 199608 138355 199613
rect 138246 199552 138294 199608
rect 138350 199552 138355 199608
rect 138246 199550 138355 199552
rect 136652 199548 136699 199550
rect 136633 199547 136699 199548
rect 138105 199547 138171 199550
rect 138289 199547 138355 199550
rect 139342 199548 139348 199612
rect 139412 199610 139418 199612
rect 139485 199610 139551 199613
rect 139412 199608 139551 199610
rect 139412 199552 139490 199608
rect 139546 199552 139551 199608
rect 139412 199550 139551 199552
rect 139412 199548 139418 199550
rect 139485 199547 139551 199550
rect 141325 199608 141391 199613
rect 141325 199552 141330 199608
rect 141386 199552 141391 199608
rect 141325 199547 141391 199552
rect 141550 199548 141556 199612
rect 141620 199610 141626 199612
rect 142705 199610 142771 199613
rect 141620 199608 142771 199610
rect 141620 199552 142710 199608
rect 142766 199552 142771 199608
rect 141620 199550 142771 199552
rect 141620 199548 141626 199550
rect 142705 199547 142771 199550
rect 147673 199610 147739 199613
rect 147814 199610 147874 199686
rect 148409 199683 148475 199686
rect 148547 199744 148613 199749
rect 148731 199748 148797 199749
rect 148547 199688 148552 199744
rect 148608 199688 148613 199744
rect 148547 199683 148613 199688
rect 148726 199684 148732 199748
rect 148796 199746 148802 199748
rect 149516 199746 149576 200094
rect 150014 200092 150020 200156
rect 150084 200154 150090 200156
rect 178309 200154 178375 200157
rect 201769 200154 201835 200157
rect 150084 200094 157626 200154
rect 150084 200092 150090 200094
rect 151302 200018 151308 200020
rect 150942 199958 151308 200018
rect 149651 199914 149717 199919
rect 149651 199884 149656 199914
rect 149712 199884 149717 199914
rect 150755 199914 150821 199919
rect 149646 199820 149652 199884
rect 149716 199882 149722 199884
rect 149927 199882 149993 199885
rect 150755 199884 150760 199914
rect 150816 199884 150821 199914
rect 150382 199882 150388 199884
rect 149716 199822 149774 199882
rect 149927 199880 150388 199882
rect 149927 199824 149932 199880
rect 149988 199824 150388 199880
rect 149927 199822 150388 199824
rect 149716 199820 149722 199822
rect 149927 199819 149993 199822
rect 150382 199820 150388 199822
rect 150452 199820 150458 199884
rect 150750 199820 150756 199884
rect 150820 199882 150826 199884
rect 150942 199882 151002 199958
rect 151302 199956 151308 199958
rect 151372 199956 151378 200020
rect 151486 199956 151492 200020
rect 151556 200018 151562 200020
rect 151556 199956 151600 200018
rect 153510 199956 153516 200020
rect 153580 200018 153586 200020
rect 153580 199958 154498 200018
rect 153580 199956 153586 199958
rect 151215 199882 151281 199885
rect 150820 199822 150878 199882
rect 150942 199880 151281 199882
rect 150942 199824 151220 199880
rect 151276 199824 151281 199880
rect 150942 199822 151281 199824
rect 150820 199820 150826 199822
rect 151215 199819 151281 199822
rect 151399 199882 151465 199885
rect 151540 199882 151600 199956
rect 152503 199916 152569 199919
rect 152276 199914 152569 199916
rect 152043 199884 152109 199885
rect 152276 199884 152508 199914
rect 152038 199882 152044 199884
rect 151399 199880 151600 199882
rect 151399 199824 151404 199880
rect 151460 199824 151600 199880
rect 151399 199822 151600 199824
rect 151952 199822 152044 199882
rect 151399 199819 151465 199822
rect 152038 199820 152044 199822
rect 152108 199820 152114 199884
rect 152222 199820 152228 199884
rect 152292 199858 152508 199884
rect 152564 199858 152569 199914
rect 152779 199914 152845 199919
rect 152779 199884 152784 199914
rect 152840 199884 152845 199914
rect 153055 199916 153121 199919
rect 153055 199914 153164 199916
rect 152292 199856 152569 199858
rect 152292 199822 152336 199856
rect 152503 199853 152569 199856
rect 152292 199820 152298 199822
rect 152774 199820 152780 199884
rect 152844 199882 152850 199884
rect 152844 199822 152902 199882
rect 153055 199858 153060 199914
rect 153116 199884 153164 199914
rect 154438 199885 154498 199958
rect 155263 199914 155329 199919
rect 153116 199858 153148 199884
rect 153055 199853 153148 199858
rect 153104 199822 153148 199853
rect 152844 199820 152850 199822
rect 153142 199820 153148 199822
rect 153212 199820 153218 199884
rect 153326 199820 153332 199884
rect 153396 199882 153402 199884
rect 153607 199882 153673 199885
rect 153396 199880 153673 199882
rect 153396 199824 153612 199880
rect 153668 199824 153673 199880
rect 153396 199822 153673 199824
rect 153396 199820 153402 199822
rect 152043 199819 152109 199820
rect 153607 199819 153673 199822
rect 153878 199820 153884 199884
rect 153948 199882 153954 199884
rect 154159 199882 154225 199885
rect 153948 199880 154225 199882
rect 153948 199824 154164 199880
rect 154220 199824 154225 199880
rect 153948 199822 154225 199824
rect 153948 199820 153954 199822
rect 154159 199819 154225 199822
rect 154435 199880 154501 199885
rect 154803 199884 154869 199885
rect 154798 199882 154804 199884
rect 154435 199824 154440 199880
rect 154496 199824 154501 199880
rect 154435 199819 154501 199824
rect 154712 199822 154804 199882
rect 154798 199820 154804 199822
rect 154868 199820 154874 199884
rect 155263 199858 155268 199914
rect 155324 199882 155329 199914
rect 157011 199914 157077 199919
rect 155534 199882 155540 199884
rect 155324 199858 155540 199882
rect 155263 199853 155540 199858
rect 155266 199822 155540 199853
rect 155534 199820 155540 199822
rect 155604 199820 155610 199884
rect 155815 199882 155881 199885
rect 156086 199882 156092 199884
rect 155815 199880 156092 199882
rect 155815 199824 155820 199880
rect 155876 199824 156092 199880
rect 155815 199822 156092 199824
rect 154803 199819 154869 199820
rect 155815 199819 155881 199822
rect 156086 199820 156092 199822
rect 156156 199820 156162 199884
rect 157011 199858 157016 199914
rect 157072 199882 157077 199914
rect 157374 199882 157380 199884
rect 157072 199858 157380 199882
rect 157011 199853 157380 199858
rect 157014 199822 157380 199853
rect 157374 199820 157380 199822
rect 157444 199820 157450 199884
rect 157566 199882 157626 200094
rect 178309 200152 201835 200154
rect 178309 200096 178314 200152
rect 178370 200096 201774 200152
rect 201830 200096 201835 200152
rect 178309 200094 201835 200096
rect 178309 200091 178375 200094
rect 201769 200091 201835 200094
rect 165286 199956 165292 200020
rect 165356 200018 165362 200020
rect 168782 200018 168788 200020
rect 165356 199958 165722 200018
rect 165356 199956 165362 199958
rect 160231 199882 160297 199885
rect 157566 199880 160297 199882
rect 157566 199824 160236 199880
rect 160292 199824 160297 199880
rect 157566 199822 160297 199824
rect 160231 199819 160297 199822
rect 160502 199820 160508 199884
rect 160572 199882 160578 199884
rect 161887 199882 161953 199885
rect 160572 199880 161953 199882
rect 160572 199824 161892 199880
rect 161948 199824 161953 199880
rect 160572 199822 161953 199824
rect 160572 199820 160578 199822
rect 161887 199819 161953 199822
rect 162342 199820 162348 199884
rect 162412 199882 162418 199884
rect 162623 199882 162689 199885
rect 163451 199884 163517 199885
rect 163446 199882 163452 199884
rect 162412 199880 162689 199882
rect 162412 199824 162628 199880
rect 162684 199824 162689 199880
rect 162412 199822 162689 199824
rect 163360 199822 163452 199882
rect 162412 199820 162418 199822
rect 162623 199819 162689 199822
rect 163446 199820 163452 199822
rect 163516 199820 163522 199884
rect 163630 199820 163636 199884
rect 163700 199882 163706 199884
rect 163819 199882 163885 199885
rect 163700 199880 163885 199882
rect 163700 199824 163824 199880
rect 163880 199824 163885 199880
rect 163700 199822 163885 199824
rect 163700 199820 163706 199822
rect 163451 199819 163517 199820
rect 163819 199819 163885 199822
rect 164366 199820 164372 199884
rect 164436 199882 164442 199884
rect 164831 199882 164897 199885
rect 165107 199884 165173 199885
rect 165102 199882 165108 199884
rect 164436 199880 164897 199882
rect 164436 199824 164836 199880
rect 164892 199824 164897 199880
rect 164436 199822 164897 199824
rect 165016 199822 165108 199882
rect 164436 199820 164442 199822
rect 164831 199819 164897 199822
rect 165102 199820 165108 199822
rect 165172 199820 165178 199884
rect 165383 199882 165449 199885
rect 165662 199882 165722 199958
rect 166398 199958 168788 200018
rect 166398 199885 166458 199958
rect 168782 199956 168788 199958
rect 168852 199956 168858 200020
rect 174670 200018 174676 200020
rect 171918 199958 174676 200018
rect 171918 199885 171978 199958
rect 174670 199956 174676 199958
rect 174740 199956 174746 200020
rect 165383 199880 165722 199882
rect 165383 199824 165388 199880
rect 165444 199824 165722 199880
rect 165383 199822 165722 199824
rect 166395 199880 166461 199885
rect 166395 199824 166400 199880
rect 166456 199824 166461 199880
rect 165107 199819 165173 199820
rect 165383 199819 165449 199822
rect 166395 199819 166461 199824
rect 166574 199820 166580 199884
rect 166644 199882 166650 199884
rect 166763 199882 166829 199885
rect 167131 199884 167197 199885
rect 167126 199882 167132 199884
rect 166644 199880 166829 199882
rect 166644 199824 166768 199880
rect 166824 199824 166829 199880
rect 166644 199822 166829 199824
rect 167040 199822 167132 199882
rect 166644 199820 166650 199822
rect 166763 199819 166829 199822
rect 167126 199820 167132 199822
rect 167196 199820 167202 199884
rect 167407 199882 167473 199885
rect 167867 199884 167933 199885
rect 167540 199882 167546 199884
rect 167407 199880 167546 199882
rect 167407 199824 167412 199880
rect 167468 199824 167546 199880
rect 167407 199822 167546 199824
rect 167131 199819 167197 199820
rect 167407 199819 167473 199822
rect 167540 199820 167546 199822
rect 167610 199820 167616 199884
rect 167862 199882 167868 199884
rect 167776 199822 167868 199882
rect 167862 199820 167868 199822
rect 167932 199820 167938 199884
rect 168966 199820 168972 199884
rect 169036 199882 169042 199884
rect 169615 199882 169681 199885
rect 169036 199880 169681 199882
rect 169036 199824 169620 199880
rect 169676 199824 169681 199880
rect 169036 199822 169681 199824
rect 169036 199820 169042 199822
rect 167867 199819 167933 199820
rect 169615 199819 169681 199822
rect 170443 199882 170509 199885
rect 170806 199882 170812 199884
rect 170443 199880 170812 199882
rect 170443 199824 170448 199880
rect 170504 199824 170812 199880
rect 170443 199822 170812 199824
rect 170443 199819 170509 199822
rect 170806 199820 170812 199822
rect 170876 199820 170882 199884
rect 171087 199882 171153 199885
rect 171547 199884 171613 199885
rect 171358 199882 171364 199884
rect 171087 199880 171364 199882
rect 171087 199824 171092 199880
rect 171148 199824 171364 199880
rect 171087 199822 171364 199824
rect 171087 199819 171153 199822
rect 171358 199820 171364 199822
rect 171428 199820 171434 199884
rect 171542 199820 171548 199884
rect 171612 199882 171618 199884
rect 171612 199822 171704 199882
rect 171915 199880 171981 199885
rect 172467 199884 172533 199885
rect 172462 199882 172468 199884
rect 171915 199824 171920 199880
rect 171976 199824 171981 199880
rect 171612 199820 171618 199822
rect 171547 199819 171613 199820
rect 171915 199819 171981 199824
rect 172376 199822 172468 199882
rect 172462 199820 172468 199822
rect 172532 199820 172538 199884
rect 172646 199820 172652 199884
rect 172716 199882 172722 199884
rect 173755 199882 173821 199885
rect 172716 199880 173821 199882
rect 172716 199824 173760 199880
rect 173816 199824 173821 199880
rect 172716 199822 173821 199824
rect 172716 199820 172722 199822
rect 172467 199819 172533 199820
rect 173755 199819 173821 199822
rect 174215 199882 174281 199885
rect 175043 199884 175109 199885
rect 175595 199884 175661 199885
rect 174486 199882 174492 199884
rect 174215 199880 174492 199882
rect 174215 199824 174220 199880
rect 174276 199824 174492 199880
rect 174215 199822 174492 199824
rect 174215 199819 174281 199822
rect 174486 199820 174492 199822
rect 174556 199820 174562 199884
rect 175038 199882 175044 199884
rect 174952 199822 175044 199882
rect 175038 199820 175044 199822
rect 175108 199820 175114 199884
rect 175590 199820 175596 199884
rect 175660 199882 175666 199884
rect 175660 199822 175752 199882
rect 175660 199820 175666 199822
rect 176326 199820 176332 199884
rect 176396 199882 176402 199884
rect 176607 199882 176673 199885
rect 176396 199880 176673 199882
rect 176396 199824 176612 199880
rect 176668 199824 176673 199880
rect 176396 199822 176673 199824
rect 176396 199820 176402 199822
rect 175043 199819 175109 199820
rect 175595 199819 175661 199820
rect 176607 199819 176673 199822
rect 176791 199882 176857 199885
rect 177849 199882 177915 199885
rect 176791 199880 177915 199882
rect 176791 199824 176796 199880
rect 176852 199824 177854 199880
rect 177910 199824 177915 199880
rect 176791 199822 177915 199824
rect 176791 199819 176857 199822
rect 177849 199819 177915 199822
rect 182766 199746 182772 199748
rect 148796 199686 148888 199746
rect 149516 199686 182772 199746
rect 148796 199684 148802 199686
rect 182766 199684 182772 199686
rect 182836 199684 182842 199748
rect 148731 199683 148797 199684
rect 147673 199608 147874 199610
rect 147673 199552 147678 199608
rect 147734 199552 147874 199608
rect 147673 199550 147874 199552
rect 148409 199610 148475 199613
rect 148550 199610 148610 199683
rect 148409 199608 148610 199610
rect 148409 199552 148414 199608
rect 148470 199552 148610 199608
rect 148409 199550 148610 199552
rect 148777 199610 148843 199613
rect 180742 199610 180748 199612
rect 148777 199608 180748 199610
rect 148777 199552 148782 199608
rect 148838 199552 180748 199608
rect 148777 199550 180748 199552
rect 147673 199547 147739 199550
rect 148409 199547 148475 199550
rect 148777 199547 148843 199550
rect 180742 199548 180748 199550
rect 180812 199548 180818 199612
rect 122598 199412 122604 199476
rect 122668 199474 122674 199476
rect 148961 199474 149027 199477
rect 149605 199476 149671 199477
rect 151721 199476 151787 199477
rect 149605 199474 149652 199476
rect 122668 199472 149027 199474
rect 122668 199416 148966 199472
rect 149022 199416 149027 199472
rect 122668 199414 149027 199416
rect 149560 199472 149652 199474
rect 149560 199416 149610 199472
rect 149560 199414 149652 199416
rect 122668 199412 122674 199414
rect 148961 199411 149027 199414
rect 149605 199412 149652 199414
rect 149716 199412 149722 199476
rect 150198 199412 150204 199476
rect 150268 199474 150274 199476
rect 151670 199474 151676 199476
rect 150268 199414 151370 199474
rect 151630 199414 151676 199474
rect 151740 199472 151787 199476
rect 151782 199416 151787 199472
rect 150268 199412 150274 199414
rect 149605 199411 149671 199412
rect 123845 199338 123911 199341
rect 150433 199338 150499 199341
rect 123845 199336 150499 199338
rect 123845 199280 123850 199336
rect 123906 199280 150438 199336
rect 150494 199280 150499 199336
rect 123845 199278 150499 199280
rect 123845 199275 123911 199278
rect 150433 199275 150499 199278
rect 123753 199202 123819 199205
rect 149881 199202 149947 199205
rect 123753 199200 149947 199202
rect 123753 199144 123758 199200
rect 123814 199144 149886 199200
rect 149942 199144 149947 199200
rect 123753 199142 149947 199144
rect 151310 199202 151370 199414
rect 151670 199412 151676 199414
rect 151740 199412 151787 199416
rect 152038 199412 152044 199476
rect 152108 199474 152114 199476
rect 154849 199474 154915 199477
rect 152108 199472 154915 199474
rect 152108 199416 154854 199472
rect 154910 199416 154915 199472
rect 152108 199414 154915 199416
rect 152108 199412 152114 199414
rect 151721 199411 151787 199412
rect 154849 199411 154915 199414
rect 156822 199412 156828 199476
rect 156892 199474 156898 199476
rect 156965 199474 157031 199477
rect 156892 199472 157031 199474
rect 156892 199416 156970 199472
rect 157026 199416 157031 199472
rect 156892 199414 157031 199416
rect 156892 199412 156898 199414
rect 156965 199411 157031 199414
rect 158897 199474 158963 199477
rect 174261 199474 174327 199477
rect 174486 199474 174492 199476
rect 158897 199472 173266 199474
rect 158897 199416 158902 199472
rect 158958 199416 173266 199472
rect 158897 199414 173266 199416
rect 158897 199411 158963 199414
rect 153878 199276 153884 199340
rect 153948 199338 153954 199340
rect 154021 199338 154087 199341
rect 153948 199336 154087 199338
rect 153948 199280 154026 199336
rect 154082 199280 154087 199336
rect 153948 199278 154087 199280
rect 153948 199276 153954 199278
rect 154021 199275 154087 199278
rect 154798 199276 154804 199340
rect 154868 199338 154874 199340
rect 154941 199338 155007 199341
rect 154868 199336 155007 199338
rect 154868 199280 154946 199336
rect 155002 199280 155007 199336
rect 154868 199278 155007 199280
rect 154868 199276 154874 199278
rect 154941 199275 155007 199278
rect 155769 199338 155835 199341
rect 156086 199338 156092 199340
rect 155769 199336 156092 199338
rect 155769 199280 155774 199336
rect 155830 199280 156092 199336
rect 155769 199278 156092 199280
rect 155769 199275 155835 199278
rect 156086 199276 156092 199278
rect 156156 199276 156162 199340
rect 157149 199338 157215 199341
rect 157374 199338 157380 199340
rect 157149 199336 157380 199338
rect 157149 199280 157154 199336
rect 157210 199280 157380 199336
rect 157149 199278 157380 199280
rect 157149 199275 157215 199278
rect 157374 199276 157380 199278
rect 157444 199276 157450 199340
rect 158294 199276 158300 199340
rect 158364 199338 158370 199340
rect 158529 199338 158595 199341
rect 158364 199336 158595 199338
rect 158364 199280 158534 199336
rect 158590 199280 158595 199336
rect 158364 199278 158595 199280
rect 158364 199276 158370 199278
rect 158529 199275 158595 199278
rect 161238 199276 161244 199340
rect 161308 199338 161314 199340
rect 162117 199338 162183 199341
rect 165153 199340 165219 199341
rect 165102 199338 165108 199340
rect 161308 199336 162183 199338
rect 161308 199280 162122 199336
rect 162178 199280 162183 199336
rect 161308 199278 162183 199280
rect 165062 199278 165108 199338
rect 165172 199336 165219 199340
rect 165214 199280 165219 199336
rect 161308 199276 161314 199278
rect 162117 199275 162183 199278
rect 165102 199276 165108 199278
rect 165172 199276 165219 199280
rect 165153 199275 165219 199276
rect 166349 199338 166415 199341
rect 170397 199340 170463 199341
rect 170857 199340 170923 199341
rect 170254 199338 170260 199340
rect 166349 199336 170260 199338
rect 166349 199280 166354 199336
rect 166410 199280 170260 199336
rect 166349 199278 170260 199280
rect 166349 199275 166415 199278
rect 170254 199276 170260 199278
rect 170324 199276 170330 199340
rect 170397 199336 170444 199340
rect 170508 199338 170514 199340
rect 170806 199338 170812 199340
rect 170397 199280 170402 199336
rect 170397 199276 170444 199280
rect 170508 199278 170554 199338
rect 170766 199278 170812 199338
rect 170876 199336 170923 199340
rect 170918 199280 170923 199336
rect 170508 199276 170514 199278
rect 170806 199276 170812 199278
rect 170876 199276 170923 199280
rect 170397 199275 170463 199276
rect 170857 199275 170923 199276
rect 171133 199338 171199 199341
rect 171358 199338 171364 199340
rect 171133 199336 171364 199338
rect 171133 199280 171138 199336
rect 171194 199280 171364 199336
rect 171133 199278 171364 199280
rect 171133 199275 171199 199278
rect 171358 199276 171364 199278
rect 171428 199276 171434 199340
rect 171726 199276 171732 199340
rect 171796 199338 171802 199340
rect 172145 199338 172211 199341
rect 171796 199336 172211 199338
rect 171796 199280 172150 199336
rect 172206 199280 172211 199336
rect 171796 199278 172211 199280
rect 171796 199276 171802 199278
rect 172145 199275 172211 199278
rect 172789 199338 172855 199341
rect 172973 199338 173039 199341
rect 172789 199336 173039 199338
rect 172789 199280 172794 199336
rect 172850 199280 172978 199336
rect 173034 199280 173039 199336
rect 172789 199278 173039 199280
rect 173206 199338 173266 199414
rect 174261 199472 174492 199474
rect 174261 199416 174266 199472
rect 174322 199416 174492 199472
rect 174261 199414 174492 199416
rect 174261 199411 174327 199414
rect 174486 199412 174492 199414
rect 174556 199412 174562 199476
rect 174670 199412 174676 199476
rect 174740 199474 174746 199476
rect 174813 199474 174879 199477
rect 174740 199472 174879 199474
rect 174740 199416 174818 199472
rect 174874 199416 174879 199472
rect 174740 199414 174879 199416
rect 174740 199412 174746 199414
rect 174813 199411 174879 199414
rect 175590 199412 175596 199476
rect 175660 199474 175666 199476
rect 176510 199474 176516 199476
rect 175660 199414 176516 199474
rect 175660 199412 175666 199414
rect 176510 199412 176516 199414
rect 176580 199412 176586 199476
rect 177297 199338 177363 199341
rect 173206 199336 177363 199338
rect 173206 199280 177302 199336
rect 177358 199280 177363 199336
rect 173206 199278 177363 199280
rect 172789 199275 172855 199278
rect 172973 199275 173039 199278
rect 177297 199275 177363 199278
rect 158253 199202 158319 199205
rect 151310 199200 158319 199202
rect 151310 199144 158258 199200
rect 158314 199144 158319 199200
rect 151310 199142 158319 199144
rect 123753 199139 123819 199142
rect 149881 199139 149947 199142
rect 158253 199139 158319 199142
rect 158529 199202 158595 199205
rect 179638 199202 179644 199204
rect 158529 199200 179644 199202
rect 158529 199144 158534 199200
rect 158590 199144 179644 199200
rect 158529 199142 179644 199144
rect 158529 199139 158595 199142
rect 179638 199140 179644 199142
rect 179708 199140 179714 199204
rect 102041 199066 102107 199069
rect 129273 199066 129339 199069
rect 102041 199064 129339 199066
rect 102041 199008 102046 199064
rect 102102 199008 129278 199064
rect 129334 199008 129339 199064
rect 102041 199006 129339 199008
rect 102041 199003 102107 199006
rect 129273 199003 129339 199006
rect 135529 199066 135595 199069
rect 136449 199068 136515 199069
rect 135846 199066 135852 199068
rect 135529 199064 135852 199066
rect 135529 199008 135534 199064
rect 135590 199008 135852 199064
rect 135529 199006 135852 199008
rect 135529 199003 135595 199006
rect 135846 199004 135852 199006
rect 135916 199004 135922 199068
rect 136398 199004 136404 199068
rect 136468 199066 136515 199068
rect 139301 199068 139367 199069
rect 139301 199066 139348 199068
rect 136468 199064 136560 199066
rect 136510 199008 136560 199064
rect 136468 199006 136560 199008
rect 139256 199064 139348 199066
rect 139256 199008 139306 199064
rect 139256 199006 139348 199008
rect 136468 199004 136515 199006
rect 136449 199003 136515 199004
rect 139301 199004 139348 199006
rect 139412 199004 139418 199068
rect 140262 199004 140268 199068
rect 140332 199066 140338 199068
rect 140681 199066 140747 199069
rect 140332 199064 140747 199066
rect 140332 199008 140686 199064
rect 140742 199008 140747 199064
rect 140332 199006 140747 199008
rect 140332 199004 140338 199006
rect 139301 199003 139367 199004
rect 140681 199003 140747 199006
rect 143441 199066 143507 199069
rect 145414 199066 145420 199068
rect 143441 199064 145420 199066
rect 143441 199008 143446 199064
rect 143502 199008 145420 199064
rect 143441 199006 145420 199008
rect 143441 199003 143507 199006
rect 145414 199004 145420 199006
rect 145484 199004 145490 199068
rect 147029 199066 147095 199069
rect 165981 199066 166047 199069
rect 166390 199066 166396 199068
rect 147029 199064 160110 199066
rect 147029 199008 147034 199064
rect 147090 199008 160110 199064
rect 147029 199006 160110 199008
rect 147029 199003 147095 199006
rect 144085 198930 144151 198933
rect 144085 198928 144194 198930
rect 144085 198872 144090 198928
rect 144146 198872 144194 198928
rect 144085 198867 144194 198872
rect 146886 198868 146892 198932
rect 146956 198930 146962 198932
rect 147213 198930 147279 198933
rect 147949 198932 148015 198933
rect 147949 198930 147996 198932
rect 146956 198928 147279 198930
rect 146956 198872 147218 198928
rect 147274 198872 147279 198928
rect 146956 198870 147279 198872
rect 147904 198928 147996 198930
rect 147904 198872 147954 198928
rect 147904 198870 147996 198872
rect 146956 198868 146962 198870
rect 147213 198867 147279 198870
rect 147949 198868 147996 198870
rect 148060 198868 148066 198932
rect 148133 198930 148199 198933
rect 148726 198930 148732 198932
rect 148133 198928 148732 198930
rect 148133 198872 148138 198928
rect 148194 198872 148732 198928
rect 148133 198870 148732 198872
rect 147949 198867 148015 198868
rect 148133 198867 148199 198870
rect 148726 198868 148732 198870
rect 148796 198868 148802 198932
rect 156873 198930 156939 198933
rect 157190 198930 157196 198932
rect 156873 198928 157196 198930
rect 156873 198872 156878 198928
rect 156934 198872 157196 198928
rect 156873 198870 157196 198872
rect 156873 198867 156939 198870
rect 157190 198868 157196 198870
rect 157260 198868 157266 198932
rect 144134 198797 144194 198867
rect 107561 198794 107627 198797
rect 136541 198794 136607 198797
rect 107561 198792 136607 198794
rect 107561 198736 107566 198792
rect 107622 198736 136546 198792
rect 136602 198736 136607 198792
rect 107561 198734 136607 198736
rect 107561 198731 107627 198734
rect 136541 198731 136607 198734
rect 139158 198732 139164 198796
rect 139228 198794 139234 198796
rect 139485 198794 139551 198797
rect 139228 198792 139551 198794
rect 139228 198736 139490 198792
rect 139546 198736 139551 198792
rect 139228 198734 139551 198736
rect 144134 198792 144243 198797
rect 144134 198736 144182 198792
rect 144238 198736 144243 198792
rect 144134 198734 144243 198736
rect 139228 198732 139234 198734
rect 139485 198731 139551 198734
rect 144177 198731 144243 198734
rect 147213 198794 147279 198797
rect 156965 198796 157031 198797
rect 150750 198794 150756 198796
rect 147213 198792 150756 198794
rect 147213 198736 147218 198792
rect 147274 198736 150756 198792
rect 147213 198734 150756 198736
rect 147213 198731 147279 198734
rect 150750 198732 150756 198734
rect 150820 198732 150826 198796
rect 156965 198792 157012 198796
rect 157076 198794 157082 198796
rect 157885 198794 157951 198797
rect 158110 198794 158116 198796
rect 156965 198736 156970 198792
rect 156965 198732 157012 198736
rect 157076 198734 157122 198794
rect 157885 198792 158116 198794
rect 157885 198736 157890 198792
rect 157946 198736 158116 198792
rect 157885 198734 158116 198736
rect 157076 198732 157082 198734
rect 156965 198731 157031 198732
rect 157885 198731 157951 198734
rect 158110 198732 158116 198734
rect 158180 198732 158186 198796
rect 160050 198794 160110 199006
rect 165981 199064 166396 199066
rect 165981 199008 165986 199064
rect 166042 199008 166396 199064
rect 165981 199006 166396 199008
rect 165981 199003 166047 199006
rect 166390 199004 166396 199006
rect 166460 199004 166466 199068
rect 172053 199066 172119 199069
rect 172697 199066 172763 199069
rect 172053 199064 172763 199066
rect 172053 199008 172058 199064
rect 172114 199008 172702 199064
rect 172758 199008 172763 199064
rect 172053 199006 172763 199008
rect 172053 199003 172119 199006
rect 172697 199003 172763 199006
rect 174445 199066 174511 199069
rect 175457 199066 175523 199069
rect 174445 199064 175523 199066
rect 174445 199008 174450 199064
rect 174506 199008 175462 199064
rect 175518 199008 175523 199064
rect 174445 199006 175523 199008
rect 174445 199003 174511 199006
rect 175457 199003 175523 199006
rect 175958 199004 175964 199068
rect 176028 199066 176034 199068
rect 176193 199066 176259 199069
rect 176469 199068 176535 199069
rect 176469 199066 176516 199068
rect 176028 199064 176259 199066
rect 176028 199008 176198 199064
rect 176254 199008 176259 199064
rect 176028 199006 176259 199008
rect 176424 199064 176516 199066
rect 176424 199008 176474 199064
rect 176424 199006 176516 199008
rect 176028 199004 176034 199006
rect 176193 199003 176259 199006
rect 176469 199004 176516 199006
rect 176580 199004 176586 199068
rect 176469 199003 176535 199004
rect 165981 198932 166047 198933
rect 165981 198930 166028 198932
rect 165936 198928 166028 198930
rect 165936 198872 165986 198928
rect 165936 198870 166028 198872
rect 165981 198868 166028 198870
rect 166092 198868 166098 198932
rect 166206 198868 166212 198932
rect 166276 198930 166282 198932
rect 166809 198930 166875 198933
rect 167821 198932 167887 198933
rect 167821 198930 167868 198932
rect 166276 198928 166875 198930
rect 166276 198872 166814 198928
rect 166870 198872 166875 198928
rect 166276 198870 166875 198872
rect 167776 198928 167868 198930
rect 167776 198872 167826 198928
rect 167776 198870 167868 198872
rect 166276 198868 166282 198870
rect 165981 198867 166047 198868
rect 166809 198867 166875 198870
rect 167821 198868 167868 198870
rect 167932 198868 167938 198932
rect 178350 198930 178356 198932
rect 170998 198870 178356 198930
rect 167821 198867 167887 198868
rect 170998 198794 171058 198870
rect 178350 198868 178356 198870
rect 178420 198868 178426 198932
rect 160050 198734 171058 198794
rect 172462 198732 172468 198796
rect 172532 198794 172538 198796
rect 173249 198794 173315 198797
rect 172532 198792 173315 198794
rect 172532 198736 173254 198792
rect 173310 198736 173315 198792
rect 172532 198734 173315 198736
rect 172532 198732 172538 198734
rect 173249 198731 173315 198734
rect 174169 198794 174235 198797
rect 199326 198794 199332 198796
rect 174169 198792 199332 198794
rect 174169 198736 174174 198792
rect 174230 198736 199332 198792
rect 174169 198734 199332 198736
rect 174169 198731 174235 198734
rect 199326 198732 199332 198734
rect 199396 198732 199402 198796
rect 133505 198660 133571 198661
rect 133454 198658 133460 198660
rect 133414 198598 133460 198658
rect 133524 198656 133571 198660
rect 139945 198658 140011 198661
rect 133566 198600 133571 198656
rect 133454 198596 133460 198598
rect 133524 198596 133571 198600
rect 133505 198595 133571 198596
rect 134014 198656 140011 198658
rect 134014 198600 139950 198656
rect 140006 198600 140011 198656
rect 134014 198598 140011 198600
rect 130878 198460 130884 198524
rect 130948 198522 130954 198524
rect 134014 198522 134074 198598
rect 139945 198595 140011 198598
rect 148910 198596 148916 198660
rect 148980 198658 148986 198660
rect 154573 198658 154639 198661
rect 148980 198656 154639 198658
rect 148980 198600 154578 198656
rect 154634 198600 154639 198656
rect 148980 198598 154639 198600
rect 148980 198596 148986 198598
rect 154573 198595 154639 198598
rect 154941 198658 155007 198661
rect 172697 198658 172763 198661
rect 186998 198658 187004 198660
rect 154941 198656 167010 198658
rect 154941 198600 154946 198656
rect 155002 198600 167010 198656
rect 154941 198598 167010 198600
rect 154941 198595 155007 198598
rect 130948 198462 134074 198522
rect 135253 198522 135319 198525
rect 144361 198522 144427 198525
rect 135253 198520 144427 198522
rect 135253 198464 135258 198520
rect 135314 198464 144366 198520
rect 144422 198464 144427 198520
rect 135253 198462 144427 198464
rect 130948 198460 130954 198462
rect 135253 198459 135319 198462
rect 144361 198459 144427 198462
rect 149421 198522 149487 198525
rect 150382 198522 150388 198524
rect 149421 198520 150388 198522
rect 149421 198464 149426 198520
rect 149482 198464 150388 198520
rect 149421 198462 150388 198464
rect 149421 198459 149487 198462
rect 150382 198460 150388 198462
rect 150452 198460 150458 198524
rect 125358 198324 125364 198388
rect 125428 198386 125434 198388
rect 145373 198386 145439 198389
rect 125428 198384 145439 198386
rect 125428 198328 145378 198384
rect 145434 198328 145439 198384
rect 125428 198326 145439 198328
rect 125428 198324 125434 198326
rect 145373 198323 145439 198326
rect 154573 198386 154639 198389
rect 161657 198386 161723 198389
rect 154573 198384 161723 198386
rect 154573 198328 154578 198384
rect 154634 198328 161662 198384
rect 161718 198328 161723 198384
rect 154573 198326 161723 198328
rect 154573 198323 154639 198326
rect 161657 198323 161723 198326
rect 125174 198188 125180 198252
rect 125244 198250 125250 198252
rect 125244 198190 138306 198250
rect 125244 198188 125250 198190
rect 124990 198052 124996 198116
rect 125060 198114 125066 198116
rect 136541 198114 136607 198117
rect 125060 198112 136607 198114
rect 125060 198056 136546 198112
rect 136602 198056 136607 198112
rect 125060 198054 136607 198056
rect 125060 198052 125066 198054
rect 136541 198051 136607 198054
rect 100569 197978 100635 197981
rect 133689 197978 133755 197981
rect 134425 197980 134491 197981
rect 134374 197978 134380 197980
rect 100569 197976 133755 197978
rect 100569 197920 100574 197976
rect 100630 197920 133694 197976
rect 133750 197920 133755 197976
rect 100569 197918 133755 197920
rect 134334 197918 134380 197978
rect 134444 197976 134491 197980
rect 134486 197920 134491 197976
rect 100569 197915 100635 197918
rect 133689 197915 133755 197918
rect 134374 197916 134380 197918
rect 134444 197916 134491 197920
rect 134558 197916 134564 197980
rect 134628 197978 134634 197980
rect 135161 197978 135227 197981
rect 134628 197976 135227 197978
rect 134628 197920 135166 197976
rect 135222 197920 135227 197976
rect 134628 197918 135227 197920
rect 134628 197916 134634 197918
rect 134425 197915 134491 197916
rect 135161 197915 135227 197918
rect 137369 197978 137435 197981
rect 137502 197978 137508 197980
rect 137369 197976 137508 197978
rect 137369 197920 137374 197976
rect 137430 197920 137508 197976
rect 137369 197918 137508 197920
rect 137369 197915 137435 197918
rect 137502 197916 137508 197918
rect 137572 197916 137578 197980
rect 133321 197842 133387 197845
rect 133638 197842 133644 197844
rect 133321 197840 133644 197842
rect 133321 197784 133326 197840
rect 133382 197784 133644 197840
rect 133321 197782 133644 197784
rect 133321 197779 133387 197782
rect 133638 197780 133644 197782
rect 133708 197780 133714 197844
rect 133873 197842 133939 197845
rect 134926 197842 134932 197844
rect 133873 197840 134932 197842
rect 133873 197784 133878 197840
rect 133934 197784 134932 197840
rect 133873 197782 134932 197784
rect 133873 197779 133939 197782
rect 134926 197780 134932 197782
rect 134996 197780 135002 197844
rect 136582 197780 136588 197844
rect 136652 197842 136658 197844
rect 137645 197842 137711 197845
rect 136652 197840 137711 197842
rect 136652 197784 137650 197840
rect 137706 197784 137711 197840
rect 136652 197782 137711 197784
rect 138246 197842 138306 198190
rect 145598 198188 145604 198252
rect 145668 198250 145674 198252
rect 157425 198250 157491 198253
rect 145668 198248 157491 198250
rect 145668 198192 157430 198248
rect 157486 198192 157491 198248
rect 145668 198190 157491 198192
rect 145668 198188 145674 198190
rect 157425 198187 157491 198190
rect 157558 198188 157564 198252
rect 157628 198250 157634 198252
rect 158253 198250 158319 198253
rect 157628 198248 158319 198250
rect 157628 198192 158258 198248
rect 158314 198192 158319 198248
rect 157628 198190 158319 198192
rect 157628 198188 157634 198190
rect 158253 198187 158319 198190
rect 139393 198116 139459 198117
rect 139342 198114 139348 198116
rect 139302 198054 139348 198114
rect 139412 198112 139459 198116
rect 139454 198056 139459 198112
rect 139342 198052 139348 198054
rect 139412 198052 139459 198056
rect 139393 198051 139459 198052
rect 139853 198114 139919 198117
rect 140078 198114 140084 198116
rect 139853 198112 140084 198114
rect 139853 198056 139858 198112
rect 139914 198056 140084 198112
rect 139853 198054 140084 198056
rect 139853 198051 139919 198054
rect 140078 198052 140084 198054
rect 140148 198052 140154 198116
rect 140313 198114 140379 198117
rect 140446 198114 140452 198116
rect 140313 198112 140452 198114
rect 140313 198056 140318 198112
rect 140374 198056 140452 198112
rect 140313 198054 140452 198056
rect 140313 198051 140379 198054
rect 140446 198052 140452 198054
rect 140516 198052 140522 198116
rect 144126 198052 144132 198116
rect 144196 198114 144202 198116
rect 156505 198114 156571 198117
rect 144196 198112 156571 198114
rect 144196 198056 156510 198112
rect 156566 198056 156571 198112
rect 144196 198054 156571 198056
rect 144196 198052 144202 198054
rect 156505 198051 156571 198054
rect 166533 198116 166599 198117
rect 166533 198112 166580 198116
rect 166644 198114 166650 198116
rect 166950 198114 167010 198598
rect 172697 198656 187004 198658
rect 172697 198600 172702 198656
rect 172758 198600 187004 198656
rect 172697 198598 187004 198600
rect 172697 198595 172763 198598
rect 186998 198596 187004 198598
rect 187068 198596 187074 198660
rect 173433 198520 173499 198525
rect 173433 198464 173438 198520
rect 173494 198464 173499 198520
rect 173433 198459 173499 198464
rect 175590 198460 175596 198524
rect 175660 198522 175666 198524
rect 176561 198522 176627 198525
rect 175660 198520 176627 198522
rect 175660 198464 176566 198520
rect 176622 198464 176627 198520
rect 175660 198462 176627 198464
rect 175660 198460 175666 198462
rect 176561 198459 176627 198462
rect 178125 198522 178191 198525
rect 187734 198522 187740 198524
rect 178125 198520 187740 198522
rect 178125 198464 178130 198520
rect 178186 198464 187740 198520
rect 178125 198462 187740 198464
rect 178125 198459 178191 198462
rect 187734 198460 187740 198462
rect 187804 198460 187810 198524
rect 169886 198188 169892 198252
rect 169956 198250 169962 198252
rect 171041 198250 171107 198253
rect 169956 198248 171107 198250
rect 169956 198192 171046 198248
rect 171102 198192 171107 198248
rect 169956 198190 171107 198192
rect 173436 198250 173496 198459
rect 174813 198386 174879 198389
rect 189390 198386 189396 198388
rect 174813 198384 189396 198386
rect 174813 198328 174818 198384
rect 174874 198328 189396 198384
rect 174813 198326 189396 198328
rect 174813 198323 174879 198326
rect 189390 198324 189396 198326
rect 189460 198324 189466 198388
rect 198958 198250 198964 198252
rect 173436 198190 198964 198250
rect 169956 198188 169962 198190
rect 171041 198187 171107 198190
rect 198958 198188 198964 198190
rect 199028 198188 199034 198252
rect 176694 198114 176700 198116
rect 166533 198056 166538 198112
rect 166533 198052 166580 198056
rect 166644 198054 166690 198114
rect 166950 198054 176700 198114
rect 166644 198052 166650 198054
rect 176694 198052 176700 198054
rect 176764 198052 176770 198116
rect 177062 198052 177068 198116
rect 177132 198114 177138 198116
rect 177389 198114 177455 198117
rect 177132 198112 177455 198114
rect 177132 198056 177394 198112
rect 177450 198056 177455 198112
rect 177132 198054 177455 198056
rect 177132 198052 177138 198054
rect 166533 198051 166599 198052
rect 177389 198051 177455 198054
rect 140998 197916 141004 197980
rect 141068 197978 141074 197980
rect 142654 197978 142660 197980
rect 141068 197918 142660 197978
rect 141068 197916 141074 197918
rect 142654 197916 142660 197918
rect 142724 197916 142730 197980
rect 144678 197916 144684 197980
rect 144748 197978 144754 197980
rect 144913 197978 144979 197981
rect 144748 197976 144979 197978
rect 144748 197920 144918 197976
rect 144974 197920 144979 197976
rect 144748 197918 144979 197920
rect 144748 197916 144754 197918
rect 144913 197915 144979 197918
rect 146753 197978 146819 197981
rect 146753 197976 167194 197978
rect 146753 197920 146758 197976
rect 146814 197920 167194 197976
rect 146753 197918 167194 197920
rect 146753 197915 146819 197918
rect 145557 197842 145623 197845
rect 138246 197840 145623 197842
rect 138246 197784 145562 197840
rect 145618 197784 145623 197840
rect 138246 197782 145623 197784
rect 136652 197780 136658 197782
rect 137645 197779 137711 197782
rect 145557 197779 145623 197782
rect 133321 197708 133387 197709
rect 133270 197644 133276 197708
rect 133340 197706 133387 197708
rect 157425 197706 157491 197709
rect 160502 197706 160508 197708
rect 133340 197704 133432 197706
rect 133382 197648 133432 197704
rect 133340 197646 133432 197648
rect 157425 197704 160508 197706
rect 157425 197648 157430 197704
rect 157486 197648 160508 197704
rect 157425 197646 160508 197648
rect 133340 197644 133387 197646
rect 133321 197643 133387 197644
rect 157425 197643 157491 197646
rect 160502 197644 160508 197646
rect 160572 197644 160578 197708
rect 167134 197706 167194 197918
rect 169150 197916 169156 197980
rect 169220 197978 169226 197980
rect 169293 197978 169359 197981
rect 169220 197976 169359 197978
rect 169220 197920 169298 197976
rect 169354 197920 169359 197976
rect 169220 197918 169359 197920
rect 169220 197916 169226 197918
rect 169293 197915 169359 197918
rect 173709 197978 173775 197981
rect 174118 197978 174124 197980
rect 173709 197976 174124 197978
rect 173709 197920 173714 197976
rect 173770 197920 174124 197976
rect 173709 197918 174124 197920
rect 173709 197915 173775 197918
rect 174118 197916 174124 197918
rect 174188 197916 174194 197980
rect 174486 197916 174492 197980
rect 174556 197978 174562 197980
rect 174997 197978 175063 197981
rect 174556 197976 175063 197978
rect 174556 197920 175002 197976
rect 175058 197920 175063 197976
rect 174556 197918 175063 197920
rect 174556 197916 174562 197918
rect 174997 197915 175063 197918
rect 176878 197916 176884 197980
rect 176948 197978 176954 197980
rect 177481 197978 177547 197981
rect 176948 197976 177547 197978
rect 176948 197920 177486 197976
rect 177542 197920 177547 197976
rect 176948 197918 177547 197920
rect 176948 197916 176954 197918
rect 177481 197915 177547 197918
rect 172881 197842 172947 197845
rect 187918 197842 187924 197844
rect 172881 197840 187924 197842
rect 172881 197784 172886 197840
rect 172942 197784 187924 197840
rect 172881 197782 187924 197784
rect 172881 197779 172947 197782
rect 187918 197780 187924 197782
rect 187988 197780 187994 197844
rect 179454 197706 179460 197708
rect 167134 197646 179460 197706
rect 179454 197644 179460 197646
rect 179524 197644 179530 197708
rect 130694 197508 130700 197572
rect 130764 197570 130770 197572
rect 143809 197570 143875 197573
rect 130764 197568 143875 197570
rect 130764 197512 143814 197568
rect 143870 197512 143875 197568
rect 130764 197510 143875 197512
rect 130764 197508 130770 197510
rect 143809 197507 143875 197510
rect 148726 197508 148732 197572
rect 148796 197570 148802 197572
rect 159173 197570 159239 197573
rect 148796 197568 159239 197570
rect 148796 197512 159178 197568
rect 159234 197512 159239 197568
rect 148796 197510 159239 197512
rect 148796 197508 148802 197510
rect 159173 197507 159239 197510
rect 162158 197508 162164 197572
rect 162228 197570 162234 197572
rect 163037 197570 163103 197573
rect 162228 197568 163103 197570
rect 162228 197512 163042 197568
rect 163098 197512 163103 197568
rect 162228 197510 163103 197512
rect 162228 197508 162234 197510
rect 163037 197507 163103 197510
rect 164550 197508 164556 197572
rect 164620 197570 164626 197572
rect 165061 197570 165127 197573
rect 164620 197568 165127 197570
rect 164620 197512 165066 197568
rect 165122 197512 165127 197568
rect 164620 197510 165127 197512
rect 164620 197508 164626 197510
rect 165061 197507 165127 197510
rect 167545 197570 167611 197573
rect 167678 197570 167684 197572
rect 167545 197568 167684 197570
rect 167545 197512 167550 197568
rect 167606 197512 167684 197568
rect 167545 197510 167684 197512
rect 167545 197507 167611 197510
rect 167678 197508 167684 197510
rect 167748 197508 167754 197572
rect 174353 197570 174419 197573
rect 174854 197570 174860 197572
rect 174353 197568 174860 197570
rect 174353 197512 174358 197568
rect 174414 197512 174860 197568
rect 174353 197510 174860 197512
rect 174353 197507 174419 197510
rect 174854 197508 174860 197510
rect 174924 197508 174930 197572
rect 176694 197508 176700 197572
rect 176764 197570 176770 197572
rect 180926 197570 180932 197572
rect 176764 197510 180932 197570
rect 176764 197508 176770 197510
rect 180926 197508 180932 197510
rect 180996 197508 181002 197572
rect 126697 197436 126763 197437
rect 126646 197434 126652 197436
rect 126606 197374 126652 197434
rect 126716 197432 126763 197436
rect 126758 197376 126763 197432
rect 126646 197372 126652 197374
rect 126716 197372 126763 197376
rect 130510 197372 130516 197436
rect 130580 197434 130586 197436
rect 135253 197434 135319 197437
rect 130580 197432 135319 197434
rect 130580 197376 135258 197432
rect 135314 197376 135319 197432
rect 130580 197374 135319 197376
rect 130580 197372 130586 197374
rect 126697 197371 126763 197372
rect 135253 197371 135319 197374
rect 153326 197372 153332 197436
rect 153396 197434 153402 197436
rect 153653 197434 153719 197437
rect 157190 197434 157196 197436
rect 153396 197432 153719 197434
rect 153396 197376 153658 197432
rect 153714 197376 153719 197432
rect 153396 197374 153719 197376
rect 153396 197372 153402 197374
rect 153653 197371 153719 197374
rect 156830 197374 157196 197434
rect 126830 197236 126836 197300
rect 126900 197298 126906 197300
rect 146477 197298 146543 197301
rect 126900 197296 146543 197298
rect 126900 197240 146482 197296
rect 146538 197240 146543 197296
rect 126900 197238 146543 197240
rect 126900 197236 126906 197238
rect 146477 197235 146543 197238
rect 156638 197236 156644 197300
rect 156708 197298 156714 197300
rect 156830 197298 156890 197374
rect 157190 197372 157196 197374
rect 157260 197372 157266 197436
rect 160870 197372 160876 197436
rect 160940 197434 160946 197436
rect 161289 197434 161355 197437
rect 160940 197432 161355 197434
rect 160940 197376 161294 197432
rect 161350 197376 161355 197432
rect 160940 197374 161355 197376
rect 160940 197372 160946 197374
rect 161289 197371 161355 197374
rect 163078 197372 163084 197436
rect 163148 197434 163154 197436
rect 163405 197434 163471 197437
rect 163148 197432 163471 197434
rect 163148 197376 163410 197432
rect 163466 197376 163471 197432
rect 163148 197374 163471 197376
rect 163148 197372 163154 197374
rect 163405 197371 163471 197374
rect 164918 197372 164924 197436
rect 164988 197434 164994 197436
rect 165245 197434 165311 197437
rect 164988 197432 165311 197434
rect 164988 197376 165250 197432
rect 165306 197376 165311 197432
rect 164988 197374 165311 197376
rect 164988 197372 164994 197374
rect 165245 197371 165311 197374
rect 168005 197436 168071 197437
rect 168005 197432 168052 197436
rect 168116 197434 168122 197436
rect 169017 197434 169083 197437
rect 169518 197434 169524 197436
rect 168005 197376 168010 197432
rect 168005 197372 168052 197376
rect 168116 197374 168162 197434
rect 169017 197432 169524 197434
rect 169017 197376 169022 197432
rect 169078 197376 169524 197432
rect 169017 197374 169524 197376
rect 168116 197372 168122 197374
rect 168005 197371 168071 197372
rect 169017 197371 169083 197374
rect 169518 197372 169524 197374
rect 169588 197372 169594 197436
rect 170070 197372 170076 197436
rect 170140 197434 170146 197436
rect 170673 197434 170739 197437
rect 170140 197432 170739 197434
rect 170140 197376 170678 197432
rect 170734 197376 170739 197432
rect 170140 197374 170739 197376
rect 170140 197372 170146 197374
rect 170673 197371 170739 197374
rect 171358 197372 171364 197436
rect 171428 197434 171434 197436
rect 171777 197434 171843 197437
rect 171428 197432 171843 197434
rect 171428 197376 171782 197432
rect 171838 197376 171843 197432
rect 171428 197374 171843 197376
rect 171428 197372 171434 197374
rect 171777 197371 171843 197374
rect 171910 197372 171916 197436
rect 171980 197434 171986 197436
rect 172329 197434 172395 197437
rect 171980 197432 172395 197434
rect 171980 197376 172334 197432
rect 172390 197376 172395 197432
rect 171980 197374 172395 197376
rect 171980 197372 171986 197374
rect 172329 197371 172395 197374
rect 172830 197372 172836 197436
rect 172900 197434 172906 197436
rect 173525 197434 173591 197437
rect 172900 197432 173591 197434
rect 172900 197376 173530 197432
rect 173586 197376 173591 197432
rect 172900 197374 173591 197376
rect 172900 197372 172906 197374
rect 173525 197371 173591 197374
rect 174302 197372 174308 197436
rect 174372 197434 174378 197436
rect 174905 197434 174971 197437
rect 174372 197432 174971 197434
rect 174372 197376 174910 197432
rect 174966 197376 174971 197432
rect 174372 197374 174971 197376
rect 174372 197372 174378 197374
rect 174905 197371 174971 197374
rect 175406 197372 175412 197436
rect 175476 197434 175482 197436
rect 176009 197434 176075 197437
rect 175476 197432 176075 197434
rect 175476 197376 176014 197432
rect 176070 197376 176075 197432
rect 175476 197374 176075 197376
rect 175476 197372 175482 197374
rect 176009 197371 176075 197374
rect 156708 197238 156890 197298
rect 161013 197300 161079 197301
rect 161013 197296 161060 197300
rect 161124 197298 161130 197300
rect 161013 197240 161018 197296
rect 156708 197236 156714 197238
rect 161013 197236 161060 197240
rect 161124 197238 161170 197298
rect 161124 197236 161130 197238
rect 163262 197236 163268 197300
rect 163332 197298 163338 197300
rect 164233 197298 164299 197301
rect 163332 197296 164299 197298
rect 163332 197240 164238 197296
rect 164294 197240 164299 197296
rect 163332 197238 164299 197240
rect 163332 197236 163338 197238
rect 161013 197235 161079 197236
rect 164233 197235 164299 197238
rect 164877 197298 164943 197301
rect 165337 197300 165403 197301
rect 165102 197298 165108 197300
rect 164877 197296 165108 197298
rect 164877 197240 164882 197296
rect 164938 197240 165108 197296
rect 164877 197238 165108 197240
rect 164877 197235 164943 197238
rect 165102 197236 165108 197238
rect 165172 197236 165178 197300
rect 165286 197236 165292 197300
rect 165356 197298 165403 197300
rect 165356 197296 165448 197298
rect 165398 197240 165448 197296
rect 165356 197238 165448 197240
rect 165356 197236 165403 197238
rect 165654 197236 165660 197300
rect 165724 197298 165730 197300
rect 166349 197298 166415 197301
rect 165724 197296 166415 197298
rect 165724 197240 166354 197296
rect 166410 197240 166415 197296
rect 165724 197238 166415 197240
rect 165724 197236 165730 197238
rect 165337 197235 165403 197236
rect 166349 197235 166415 197238
rect 167310 197236 167316 197300
rect 167380 197298 167386 197300
rect 168281 197298 168347 197301
rect 167380 197296 168347 197298
rect 167380 197240 168286 197296
rect 168342 197240 168347 197296
rect 167380 197238 168347 197240
rect 167380 197236 167386 197238
rect 168281 197235 168347 197238
rect 169334 197236 169340 197300
rect 169404 197298 169410 197300
rect 169569 197298 169635 197301
rect 170397 197300 170463 197301
rect 172973 197300 173039 197301
rect 170397 197298 170444 197300
rect 169404 197296 169635 197298
rect 169404 197240 169574 197296
rect 169630 197240 169635 197296
rect 169404 197238 169635 197240
rect 170352 197296 170444 197298
rect 170352 197240 170402 197296
rect 170352 197238 170444 197240
rect 169404 197236 169410 197238
rect 169569 197235 169635 197238
rect 170397 197236 170444 197238
rect 170508 197236 170514 197300
rect 172973 197298 173020 197300
rect 172928 197296 173020 197298
rect 172928 197240 172978 197296
rect 172928 197238 173020 197240
rect 172973 197236 173020 197238
rect 173084 197236 173090 197300
rect 173157 197298 173223 197301
rect 174997 197300 175063 197301
rect 173382 197298 173388 197300
rect 173157 197296 173388 197298
rect 173157 197240 173162 197296
rect 173218 197240 173388 197296
rect 173157 197238 173388 197240
rect 170397 197235 170463 197236
rect 172973 197235 173039 197236
rect 173157 197235 173223 197238
rect 173382 197236 173388 197238
rect 173452 197236 173458 197300
rect 174997 197298 175044 197300
rect 174952 197296 175044 197298
rect 174952 197240 175002 197296
rect 174952 197238 175044 197240
rect 174997 197236 175044 197238
rect 175108 197236 175114 197300
rect 175457 197298 175523 197301
rect 175774 197298 175780 197300
rect 175457 197296 175780 197298
rect 175457 197240 175462 197296
rect 175518 197240 175780 197296
rect 175457 197238 175780 197240
rect 174997 197235 175063 197236
rect 175457 197235 175523 197238
rect 175774 197236 175780 197238
rect 175844 197236 175850 197300
rect 130469 197162 130535 197165
rect 151997 197162 152063 197165
rect 130469 197160 152063 197162
rect 130469 197104 130474 197160
rect 130530 197104 152002 197160
rect 152058 197104 152063 197160
rect 130469 197102 152063 197104
rect 130469 197099 130535 197102
rect 151997 197099 152063 197102
rect 160502 197100 160508 197164
rect 160572 197162 160578 197164
rect 168189 197162 168255 197165
rect 160572 197160 168255 197162
rect 160572 197104 168194 197160
rect 168250 197104 168255 197160
rect 160572 197102 168255 197104
rect 160572 197100 160578 197102
rect 168189 197099 168255 197102
rect 176745 197162 176811 197165
rect 193254 197162 193260 197164
rect 176745 197160 193260 197162
rect 176745 197104 176750 197160
rect 176806 197104 193260 197160
rect 176745 197102 193260 197104
rect 176745 197099 176811 197102
rect 193254 197100 193260 197102
rect 193324 197100 193330 197164
rect 104249 197026 104315 197029
rect 134517 197026 134583 197029
rect 104249 197024 134583 197026
rect 104249 196968 104254 197024
rect 104310 196968 134522 197024
rect 134578 196968 134583 197024
rect 104249 196966 134583 196968
rect 104249 196963 104315 196966
rect 134517 196963 134583 196966
rect 140814 196964 140820 197028
rect 140884 197026 140890 197028
rect 143574 197026 143580 197028
rect 140884 196966 143580 197026
rect 140884 196964 140890 196966
rect 143574 196964 143580 196966
rect 143644 196964 143650 197028
rect 149830 196964 149836 197028
rect 149900 197026 149906 197028
rect 150065 197026 150131 197029
rect 149900 197024 150131 197026
rect 149900 196968 150070 197024
rect 150126 196968 150131 197024
rect 149900 196966 150131 196968
rect 149900 196964 149906 196966
rect 150065 196963 150131 196966
rect 151302 196964 151308 197028
rect 151372 197026 151378 197028
rect 178166 197026 178172 197028
rect 151372 196966 178172 197026
rect 151372 196964 151378 196966
rect 178166 196964 178172 196966
rect 178236 196964 178242 197028
rect 107469 196890 107535 196893
rect 138565 196890 138631 196893
rect 107469 196888 138631 196890
rect 107469 196832 107474 196888
rect 107530 196832 138570 196888
rect 138626 196832 138631 196888
rect 107469 196830 138631 196832
rect 107469 196827 107535 196830
rect 138565 196827 138631 196830
rect 149462 196828 149468 196892
rect 149532 196890 149538 196892
rect 157517 196890 157583 196893
rect 149532 196888 157583 196890
rect 149532 196832 157522 196888
rect 157578 196832 157583 196888
rect 149532 196830 157583 196832
rect 149532 196828 149538 196830
rect 157517 196827 157583 196830
rect 164969 196890 165035 196893
rect 198733 196890 198799 196893
rect 164969 196888 198799 196890
rect 164969 196832 164974 196888
rect 165030 196832 198738 196888
rect 198794 196832 198799 196888
rect 164969 196830 198799 196832
rect 164969 196827 165035 196830
rect 198733 196827 198799 196830
rect 118601 196754 118667 196757
rect 151670 196754 151676 196756
rect 118601 196752 151676 196754
rect 118601 196696 118606 196752
rect 118662 196696 151676 196752
rect 118601 196694 151676 196696
rect 118601 196691 118667 196694
rect 151670 196692 151676 196694
rect 151740 196692 151746 196756
rect 157701 196754 157767 196757
rect 157926 196754 157932 196756
rect 157701 196752 157932 196754
rect 157701 196696 157706 196752
rect 157762 196696 157932 196752
rect 157701 196694 157932 196696
rect 157701 196691 157767 196694
rect 157926 196692 157932 196694
rect 157996 196692 158002 196756
rect 158846 196692 158852 196756
rect 158916 196754 158922 196756
rect 159725 196754 159791 196757
rect 158916 196752 159791 196754
rect 158916 196696 159730 196752
rect 159786 196696 159791 196752
rect 158916 196694 159791 196696
rect 158916 196692 158922 196694
rect 159725 196691 159791 196694
rect 161974 196692 161980 196756
rect 162044 196754 162050 196756
rect 162485 196754 162551 196757
rect 162044 196752 162551 196754
rect 162044 196696 162490 196752
rect 162546 196696 162551 196752
rect 162044 196694 162551 196696
rect 162044 196692 162050 196694
rect 162485 196691 162551 196694
rect 166901 196754 166967 196757
rect 200113 196754 200179 196757
rect 166901 196752 200179 196754
rect 166901 196696 166906 196752
rect 166962 196696 200118 196752
rect 200174 196696 200179 196752
rect 166901 196694 200179 196696
rect 166901 196691 166967 196694
rect 200113 196691 200179 196694
rect 118550 196556 118556 196620
rect 118620 196618 118626 196620
rect 152641 196618 152707 196621
rect 118620 196616 152707 196618
rect 118620 196560 152646 196616
rect 152702 196560 152707 196616
rect 118620 196558 152707 196560
rect 118620 196556 118626 196558
rect 152641 196555 152707 196558
rect 159030 196556 159036 196620
rect 159100 196618 159106 196620
rect 159449 196618 159515 196621
rect 159100 196616 159515 196618
rect 159100 196560 159454 196616
rect 159510 196560 159515 196616
rect 159100 196558 159515 196560
rect 159100 196556 159106 196558
rect 159449 196555 159515 196558
rect 168782 196556 168788 196620
rect 168852 196618 168858 196620
rect 200205 196618 200271 196621
rect 168852 196616 200271 196618
rect 168852 196560 200210 196616
rect 200266 196560 200271 196616
rect 168852 196558 200271 196560
rect 168852 196556 168858 196558
rect 200205 196555 200271 196558
rect 128997 196482 129063 196485
rect 142470 196482 142476 196484
rect 128997 196480 142476 196482
rect 128997 196424 129002 196480
rect 129058 196424 142476 196480
rect 128997 196422 142476 196424
rect 128997 196419 129063 196422
rect 142470 196420 142476 196422
rect 142540 196420 142546 196484
rect 149646 196420 149652 196484
rect 149716 196482 149722 196484
rect 149789 196482 149855 196485
rect 149716 196480 149855 196482
rect 149716 196424 149794 196480
rect 149850 196424 149855 196480
rect 149716 196422 149855 196424
rect 149716 196420 149722 196422
rect 149789 196419 149855 196422
rect 132677 196210 132743 196213
rect 133086 196210 133092 196212
rect 132677 196208 133092 196210
rect 132677 196152 132682 196208
rect 132738 196152 133092 196208
rect 132677 196150 133092 196152
rect 132677 196147 132743 196150
rect 133086 196148 133092 196150
rect 133156 196148 133162 196212
rect 131614 196012 131620 196076
rect 131684 196074 131690 196076
rect 132401 196074 132467 196077
rect 131684 196072 132467 196074
rect 131684 196016 132406 196072
rect 132462 196016 132467 196072
rect 131684 196014 132467 196016
rect 131684 196012 131690 196014
rect 132401 196011 132467 196014
rect 132861 196074 132927 196077
rect 133270 196074 133276 196076
rect 132861 196072 133276 196074
rect 132861 196016 132866 196072
rect 132922 196016 133276 196072
rect 132861 196014 133276 196016
rect 132861 196011 132927 196014
rect 133270 196012 133276 196014
rect 133340 196012 133346 196076
rect 140814 196012 140820 196076
rect 140884 196074 140890 196076
rect 141969 196074 142035 196077
rect 140884 196072 142035 196074
rect 140884 196016 141974 196072
rect 142030 196016 142035 196072
rect 140884 196014 142035 196016
rect 140884 196012 140890 196014
rect 141969 196011 142035 196014
rect 145230 196012 145236 196076
rect 145300 196074 145306 196076
rect 147806 196074 147812 196076
rect 145300 196014 147812 196074
rect 145300 196012 145306 196014
rect 147806 196012 147812 196014
rect 147876 196012 147882 196076
rect 151261 196074 151327 196077
rect 151486 196074 151492 196076
rect 151261 196072 151492 196074
rect 151261 196016 151266 196072
rect 151322 196016 151492 196072
rect 151261 196014 151492 196016
rect 151261 196011 151327 196014
rect 151486 196012 151492 196014
rect 151556 196012 151562 196076
rect 131798 195876 131804 195940
rect 131868 195938 131874 195940
rect 148542 195938 148548 195940
rect 131868 195878 148548 195938
rect 131868 195876 131874 195878
rect 148542 195876 148548 195878
rect 148612 195876 148618 195940
rect 176837 195938 176903 195941
rect 198774 195938 198780 195940
rect 176837 195936 198780 195938
rect 176837 195880 176842 195936
rect 176898 195880 198780 195936
rect 176837 195878 198780 195880
rect 176837 195875 176903 195878
rect 198774 195876 198780 195878
rect 198844 195876 198850 195940
rect 128118 195740 128124 195804
rect 128188 195802 128194 195804
rect 146845 195802 146911 195805
rect 128188 195800 146911 195802
rect 128188 195744 146850 195800
rect 146906 195744 146911 195800
rect 128188 195742 146911 195744
rect 128188 195740 128194 195742
rect 146845 195739 146911 195742
rect 175089 195802 175155 195805
rect 197302 195802 197308 195804
rect 175089 195800 197308 195802
rect 175089 195744 175094 195800
rect 175150 195744 197308 195800
rect 175089 195742 197308 195744
rect 175089 195739 175155 195742
rect 197302 195740 197308 195742
rect 197372 195740 197378 195804
rect 132166 195604 132172 195668
rect 132236 195666 132242 195668
rect 150341 195666 150407 195669
rect 132236 195664 150407 195666
rect 132236 195608 150346 195664
rect 150402 195608 150407 195664
rect 132236 195606 150407 195608
rect 132236 195604 132242 195606
rect 150341 195603 150407 195606
rect 150801 195666 150867 195669
rect 151118 195666 151124 195668
rect 150801 195664 151124 195666
rect 150801 195608 150806 195664
rect 150862 195608 151124 195664
rect 150801 195606 151124 195608
rect 150801 195603 150867 195606
rect 151118 195604 151124 195606
rect 151188 195604 151194 195668
rect 156270 195604 156276 195668
rect 156340 195666 156346 195668
rect 158805 195666 158871 195669
rect 156340 195664 158871 195666
rect 156340 195608 158810 195664
rect 158866 195608 158871 195664
rect 156340 195606 158871 195608
rect 156340 195604 156346 195606
rect 158805 195603 158871 195606
rect 176285 195666 176351 195669
rect 200614 195666 200620 195668
rect 176285 195664 200620 195666
rect 176285 195608 176290 195664
rect 176346 195608 200620 195664
rect 176285 195606 200620 195608
rect 176285 195603 176351 195606
rect 200614 195604 200620 195606
rect 200684 195604 200690 195668
rect 126462 195468 126468 195532
rect 126532 195530 126538 195532
rect 146109 195530 146175 195533
rect 126532 195528 146175 195530
rect 126532 195472 146114 195528
rect 146170 195472 146175 195528
rect 126532 195470 146175 195472
rect 126532 195468 126538 195470
rect 146109 195467 146175 195470
rect 147254 195468 147260 195532
rect 147324 195530 147330 195532
rect 160185 195530 160251 195533
rect 147324 195528 160251 195530
rect 147324 195472 160190 195528
rect 160246 195472 160251 195528
rect 147324 195470 160251 195472
rect 147324 195468 147330 195470
rect 160185 195467 160251 195470
rect 176326 195468 176332 195532
rect 176396 195530 176402 195532
rect 200982 195530 200988 195532
rect 176396 195470 200988 195530
rect 176396 195468 176402 195470
rect 200982 195468 200988 195470
rect 201052 195468 201058 195532
rect 114277 195394 114343 195397
rect 128721 195394 128787 195397
rect 114277 195392 128787 195394
rect 114277 195336 114282 195392
rect 114338 195336 128726 195392
rect 128782 195336 128787 195392
rect 114277 195334 128787 195336
rect 114277 195331 114343 195334
rect 128721 195331 128787 195334
rect 141969 195394 142035 195397
rect 142838 195394 142844 195396
rect 141969 195392 142844 195394
rect 141969 195336 141974 195392
rect 142030 195336 142844 195392
rect 141969 195334 142844 195336
rect 141969 195331 142035 195334
rect 142838 195332 142844 195334
rect 142908 195332 142914 195396
rect 144085 195394 144151 195397
rect 144678 195394 144684 195396
rect 144085 195392 144684 195394
rect 144085 195336 144090 195392
rect 144146 195336 144684 195392
rect 144085 195334 144684 195336
rect 144085 195331 144151 195334
rect 144678 195332 144684 195334
rect 144748 195332 144754 195396
rect 154849 195394 154915 195397
rect 182582 195394 182588 195396
rect 154849 195392 182588 195394
rect 154849 195336 154854 195392
rect 154910 195336 182588 195392
rect 154849 195334 182588 195336
rect 154849 195331 154915 195334
rect 182582 195332 182588 195334
rect 182652 195332 182658 195396
rect 124070 195196 124076 195260
rect 124140 195258 124146 195260
rect 157333 195258 157399 195261
rect 124140 195256 157399 195258
rect 124140 195200 157338 195256
rect 157394 195200 157399 195256
rect 124140 195198 157399 195200
rect 124140 195196 124146 195198
rect 157333 195195 157399 195198
rect 175181 195258 175247 195261
rect 200798 195258 200804 195260
rect 175181 195256 200804 195258
rect 175181 195200 175186 195256
rect 175242 195200 200804 195256
rect 175181 195198 200804 195200
rect 175181 195195 175247 195198
rect 200798 195196 200804 195198
rect 200868 195196 200874 195260
rect 137093 195122 137159 195125
rect 141969 195122 142035 195125
rect 137093 195120 142035 195122
rect 137093 195064 137098 195120
rect 137154 195064 141974 195120
rect 142030 195064 142035 195120
rect 137093 195062 142035 195064
rect 137093 195059 137159 195062
rect 141969 195059 142035 195062
rect 177113 195122 177179 195125
rect 196014 195122 196020 195124
rect 177113 195120 196020 195122
rect 177113 195064 177118 195120
rect 177174 195064 196020 195120
rect 177113 195062 196020 195064
rect 177113 195059 177179 195062
rect 196014 195060 196020 195062
rect 196084 195060 196090 195124
rect 124806 194108 124812 194172
rect 124876 194170 124882 194172
rect 143533 194170 143599 194173
rect 124876 194168 143599 194170
rect 124876 194112 143538 194168
rect 143594 194112 143599 194168
rect 124876 194110 143599 194112
rect 124876 194108 124882 194110
rect 143533 194107 143599 194110
rect 130326 193972 130332 194036
rect 130396 194034 130402 194036
rect 149513 194034 149579 194037
rect 130396 194032 149579 194034
rect 130396 193976 149518 194032
rect 149574 193976 149579 194032
rect 130396 193974 149579 193976
rect 130396 193972 130402 193974
rect 149513 193971 149579 193974
rect 155033 194034 155099 194037
rect 155718 194034 155724 194036
rect 155033 194032 155724 194034
rect 155033 193976 155038 194032
rect 155094 193976 155724 194032
rect 155033 193974 155724 193976
rect 155033 193971 155099 193974
rect 155718 193972 155724 193974
rect 155788 193972 155794 194036
rect 168557 194034 168623 194037
rect 201718 194034 201724 194036
rect 168557 194032 201724 194034
rect 168557 193976 168562 194032
rect 168618 193976 201724 194032
rect 168557 193974 201724 193976
rect 168557 193971 168623 193974
rect 201718 193972 201724 193974
rect 201788 193972 201794 194036
rect 104709 193898 104775 193901
rect 128077 193898 128143 193901
rect 104709 193896 128143 193898
rect 104709 193840 104714 193896
rect 104770 193840 128082 193896
rect 128138 193840 128143 193896
rect 104709 193838 128143 193840
rect 104709 193835 104775 193838
rect 128077 193835 128143 193838
rect 167913 193898 167979 193901
rect 201534 193898 201540 193900
rect 167913 193896 201540 193898
rect 167913 193840 167918 193896
rect 167974 193840 201540 193896
rect 167913 193838 201540 193840
rect 167913 193835 167979 193838
rect 201534 193836 201540 193838
rect 201604 193836 201610 193900
rect 143993 193218 144059 193221
rect 144494 193218 144500 193220
rect 143993 193216 144500 193218
rect 143993 193160 143998 193216
rect 144054 193160 144500 193216
rect 143993 193158 144500 193160
rect 143993 193155 144059 193158
rect 144494 193156 144500 193158
rect 144564 193156 144570 193220
rect 167126 193156 167132 193220
rect 167196 193218 167202 193220
rect 179689 193218 179755 193221
rect 167196 193216 179755 193218
rect 167196 193160 179694 193216
rect 179750 193160 179755 193216
rect 167196 193158 179755 193160
rect 167196 193156 167202 193158
rect 179689 193155 179755 193158
rect 177757 193082 177823 193085
rect 205725 193082 205791 193085
rect 177757 193080 205791 193082
rect 177757 193024 177762 193080
rect 177818 193024 205730 193080
rect 205786 193024 205791 193080
rect 177757 193022 205791 193024
rect 177757 193019 177823 193022
rect 205725 193019 205791 193022
rect 177021 192946 177087 192949
rect 205909 192946 205975 192949
rect 177021 192944 205975 192946
rect 177021 192888 177026 192944
rect 177082 192888 205914 192944
rect 205970 192888 205975 192944
rect 177021 192886 205975 192888
rect 177021 192883 177087 192886
rect 205909 192883 205975 192886
rect 112345 192810 112411 192813
rect 141601 192810 141667 192813
rect 112345 192808 141667 192810
rect 112345 192752 112350 192808
rect 112406 192752 141606 192808
rect 141662 192752 141667 192808
rect 112345 192750 141667 192752
rect 112345 192747 112411 192750
rect 141601 192747 141667 192750
rect 176561 192810 176627 192813
rect 206001 192810 206067 192813
rect 176561 192808 206067 192810
rect 176561 192752 176566 192808
rect 176622 192752 206006 192808
rect 206062 192752 206067 192808
rect 176561 192750 206067 192752
rect 176561 192747 176627 192750
rect 206001 192747 206067 192750
rect 111333 192674 111399 192677
rect 141325 192674 141391 192677
rect 111333 192672 141391 192674
rect 111333 192616 111338 192672
rect 111394 192616 141330 192672
rect 141386 192616 141391 192672
rect 111333 192614 141391 192616
rect 111333 192611 111399 192614
rect 141325 192611 141391 192614
rect 173157 192674 173223 192677
rect 204253 192674 204319 192677
rect 173157 192672 204319 192674
rect 173157 192616 173162 192672
rect 173218 192616 204258 192672
rect 204314 192616 204319 192672
rect 173157 192614 204319 192616
rect 173157 192611 173223 192614
rect 204253 192611 204319 192614
rect 108297 192538 108363 192541
rect 142797 192538 142863 192541
rect 108297 192536 142863 192538
rect 108297 192480 108302 192536
rect 108358 192480 142802 192536
rect 142858 192480 142863 192536
rect 108297 192478 142863 192480
rect 108297 192475 108363 192478
rect 142797 192475 142863 192478
rect 174353 192538 174419 192541
rect 205817 192538 205883 192541
rect 174353 192536 205883 192538
rect 174353 192480 174358 192536
rect 174414 192480 205822 192536
rect 205878 192480 205883 192536
rect 174353 192478 205883 192480
rect 174353 192475 174419 192478
rect 205817 192475 205883 192478
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 153694 191252 153700 191316
rect 153764 191314 153770 191316
rect 154021 191314 154087 191317
rect 153764 191312 154087 191314
rect 153764 191256 154026 191312
rect 154082 191256 154087 191312
rect 153764 191254 154087 191256
rect 153764 191252 153770 191254
rect 154021 191251 154087 191254
rect 135713 191178 135779 191181
rect 136214 191178 136220 191180
rect 135713 191176 136220 191178
rect 135713 191120 135718 191176
rect 135774 191120 136220 191176
rect 135713 191118 136220 191120
rect 135713 191115 135779 191118
rect 136214 191116 136220 191118
rect 136284 191116 136290 191180
rect 148174 191116 148180 191180
rect 148244 191178 148250 191180
rect 148593 191178 148659 191181
rect 148244 191176 148659 191178
rect 148244 191120 148598 191176
rect 148654 191120 148659 191176
rect 148244 191118 148659 191120
rect 148244 191116 148250 191118
rect 148593 191115 148659 191118
rect 162945 191178 163011 191181
rect 163446 191178 163452 191180
rect 162945 191176 163452 191178
rect 162945 191120 162950 191176
rect 163006 191120 163452 191176
rect 162945 191118 163452 191120
rect 162945 191115 163011 191118
rect 163446 191116 163452 191118
rect 163516 191116 163522 191180
rect 164233 191178 164299 191181
rect 164693 191180 164759 191181
rect 164366 191178 164372 191180
rect 164233 191176 164372 191178
rect 164233 191120 164238 191176
rect 164294 191120 164372 191176
rect 164233 191118 164372 191120
rect 164233 191115 164299 191118
rect 164366 191116 164372 191118
rect 164436 191116 164442 191180
rect 164693 191176 164740 191180
rect 164804 191178 164810 191180
rect 164693 191120 164698 191176
rect 164693 191116 164740 191120
rect 164804 191118 164850 191178
rect 164804 191116 164810 191118
rect 164693 191115 164759 191116
rect 135478 190980 135484 191044
rect 135548 191042 135554 191044
rect 135989 191042 136055 191045
rect 135548 191040 136055 191042
rect 135548 190984 135994 191040
rect 136050 190984 136055 191040
rect 135548 190982 136055 190984
rect 135548 190980 135554 190982
rect 135989 190979 136055 190982
rect 148358 190980 148364 191044
rect 148428 191042 148434 191044
rect 149053 191042 149119 191045
rect 148428 191040 149119 191042
rect 148428 190984 149058 191040
rect 149114 190984 149119 191040
rect 148428 190982 149119 190984
rect 148428 190980 148434 190982
rect 149053 190979 149119 190982
rect 153653 190906 153719 190909
rect 154062 190906 154068 190908
rect 153653 190904 154068 190906
rect 153653 190848 153658 190904
rect 153714 190848 154068 190904
rect 153653 190846 154068 190848
rect 153653 190843 153719 190846
rect 154062 190844 154068 190846
rect 154132 190844 154138 190908
rect 160502 190572 160508 190636
rect 160572 190634 160578 190636
rect 161238 190634 161244 190636
rect 160572 190574 161244 190634
rect 160572 190572 160578 190574
rect 161238 190572 161244 190574
rect 161308 190572 161314 190636
rect 160737 190500 160803 190501
rect 160686 190498 160692 190500
rect 160646 190438 160692 190498
rect 160756 190496 160803 190500
rect 160798 190440 160803 190496
rect 160686 190436 160692 190438
rect 160756 190436 160803 190440
rect 160737 190435 160803 190436
rect 161381 190362 161447 190365
rect 161336 190360 161490 190362
rect 161336 190304 161386 190360
rect 161442 190304 161490 190360
rect 161336 190302 161490 190304
rect 161381 190299 161490 190302
rect 161430 190228 161490 190299
rect 161422 190164 161428 190228
rect 161492 190164 161498 190228
rect 110965 189682 111031 189685
rect 143574 189682 143580 189684
rect 110965 189680 143580 189682
rect 110965 189624 110970 189680
rect 111026 189624 143580 189680
rect 110965 189622 143580 189624
rect 110965 189619 111031 189622
rect 143574 189620 143580 189622
rect 143644 189620 143650 189684
rect 153837 189412 153903 189413
rect 153837 189408 153884 189412
rect 153948 189410 153954 189412
rect 163589 189410 163655 189413
rect 163998 189410 164004 189412
rect 153837 189352 153842 189408
rect 153837 189348 153884 189352
rect 153948 189350 153994 189410
rect 163589 189408 164004 189410
rect 163589 189352 163594 189408
rect 163650 189352 164004 189408
rect 163589 189350 164004 189352
rect 153948 189348 153954 189350
rect 153837 189347 153903 189348
rect 163589 189347 163655 189350
rect 163998 189348 164004 189350
rect 164068 189348 164074 189412
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 140998 188804 141004 188868
rect 141068 188866 141074 188868
rect 141785 188866 141851 188869
rect 141068 188864 141851 188866
rect 141068 188808 141790 188864
rect 141846 188808 141851 188864
rect 141068 188806 141851 188808
rect 141068 188804 141074 188806
rect 141785 188803 141851 188806
rect 152181 183562 152247 183565
rect 152406 183562 152412 183564
rect 152181 183560 152412 183562
rect 152181 183504 152186 183560
rect 152242 183504 152412 183560
rect 152181 183502 152412 183504
rect 152181 183499 152247 183502
rect 152406 183500 152412 183502
rect 152476 183500 152482 183564
rect 138749 183290 138815 183293
rect 138974 183290 138980 183292
rect 138749 183288 138980 183290
rect 138749 183232 138754 183288
rect 138810 183232 138980 183288
rect 138749 183230 138980 183232
rect 138749 183227 138815 183230
rect 138974 183228 138980 183230
rect 139044 183228 139050 183292
rect 161381 180844 161447 180845
rect 161381 180842 161428 180844
rect 161336 180840 161428 180842
rect 161492 180842 161498 180844
rect 161336 180784 161386 180840
rect 161336 180782 161428 180784
rect 161381 180780 161428 180782
rect 161492 180782 161574 180842
rect 161492 180780 161498 180782
rect 161381 180779 161447 180780
rect 161381 180706 161447 180709
rect 161336 180704 161490 180706
rect 161336 180648 161386 180704
rect 161442 180648 161490 180704
rect 161336 180646 161490 180648
rect 161381 180643 161490 180646
rect 161430 180572 161490 180643
rect 161422 180508 161428 180572
rect 161492 180508 161498 180572
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 161381 171188 161447 171189
rect 161381 171186 161428 171188
rect 161336 171184 161428 171186
rect 161492 171186 161498 171188
rect 161336 171128 161386 171184
rect 161336 171126 161428 171128
rect 161381 171124 161428 171126
rect 161492 171126 161574 171186
rect 161492 171124 161498 171126
rect 161381 171123 161447 171124
rect 161381 171050 161447 171053
rect 161336 171048 161490 171050
rect 161336 170992 161386 171048
rect 161442 170992 161490 171048
rect 161336 170990 161490 170992
rect 161381 170987 161490 170990
rect 161430 170916 161490 170987
rect 161422 170852 161428 170916
rect 161492 170852 161498 170916
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 161381 161532 161447 161533
rect 161381 161530 161428 161532
rect 161336 161528 161428 161530
rect 161492 161530 161498 161532
rect 161336 161472 161386 161528
rect 161336 161470 161428 161472
rect 161381 161468 161428 161470
rect 161492 161470 161574 161530
rect 161492 161468 161498 161470
rect 161381 161467 161447 161468
rect 161381 161394 161447 161397
rect 161336 161392 161490 161394
rect 161336 161336 161386 161392
rect 161442 161336 161490 161392
rect 161336 161334 161490 161336
rect 161381 161331 161490 161334
rect 161430 161260 161490 161331
rect 161422 161196 161428 161260
rect 161492 161196 161498 161260
rect 164601 152690 164667 152693
rect 186078 152690 186084 152692
rect 164601 152688 186084 152690
rect 164601 152632 164606 152688
rect 164662 152632 186084 152688
rect 164601 152630 186084 152632
rect 164601 152627 164667 152630
rect 186078 152628 186084 152630
rect 186148 152628 186154 152692
rect 580349 152690 580415 152693
rect 583520 152690 584960 152780
rect 580349 152688 584960 152690
rect 580349 152632 580354 152688
rect 580410 152632 584960 152688
rect 580349 152630 584960 152632
rect 580349 152627 580415 152630
rect 163129 152554 163195 152557
rect 185158 152554 185164 152556
rect 163129 152552 185164 152554
rect 163129 152496 163134 152552
rect 163190 152496 185164 152552
rect 163129 152494 185164 152496
rect 163129 152491 163195 152494
rect 185158 152492 185164 152494
rect 185228 152492 185234 152556
rect 583520 152540 584960 152630
rect 161657 152418 161723 152421
rect 185342 152418 185348 152420
rect 161657 152416 185348 152418
rect 161657 152360 161662 152416
rect 161718 152360 185348 152416
rect 161657 152358 185348 152360
rect 161657 152355 161723 152358
rect 185342 152356 185348 152358
rect 185412 152356 185418 152420
rect 161381 151876 161447 151877
rect 161381 151874 161428 151876
rect 161336 151872 161428 151874
rect 161492 151874 161498 151876
rect 161336 151816 161386 151872
rect 161336 151814 161428 151816
rect 161381 151812 161428 151814
rect 161492 151814 161574 151874
rect 161492 151812 161498 151814
rect 161381 151811 161447 151812
rect 161381 151738 161447 151741
rect 161336 151736 161490 151738
rect 161336 151680 161386 151736
rect 161442 151680 161490 151736
rect 161336 151678 161490 151680
rect 161381 151675 161490 151678
rect 161430 151604 161490 151675
rect 161422 151540 161428 151604
rect 161492 151540 161498 151604
rect 179137 150378 179203 150381
rect 203006 150378 203012 150380
rect 179137 150376 203012 150378
rect 179137 150320 179142 150376
rect 179198 150320 203012 150376
rect 179137 150318 203012 150320
rect 179137 150315 179203 150318
rect 203006 150316 203012 150318
rect 203076 150316 203082 150380
rect 158529 150242 158595 150245
rect 182950 150242 182956 150244
rect 158529 150240 182956 150242
rect 158529 150184 158534 150240
rect 158590 150184 182956 150240
rect 158529 150182 182956 150184
rect 158529 150179 158595 150182
rect 182950 150180 182956 150182
rect 183020 150180 183026 150244
rect 155033 150106 155099 150109
rect 181110 150106 181116 150108
rect 155033 150104 181116 150106
rect 155033 150048 155038 150104
rect 155094 150048 181116 150104
rect 155033 150046 181116 150048
rect 155033 150043 155099 150046
rect 181110 150044 181116 150046
rect 181180 150044 181186 150108
rect 157149 149970 157215 149973
rect 183134 149970 183140 149972
rect 157149 149968 183140 149970
rect -960 149834 480 149924
rect 157149 149912 157154 149968
rect 157210 149912 183140 149968
rect 157149 149910 183140 149912
rect 157149 149907 157215 149910
rect 183134 149908 183140 149910
rect 183204 149908 183210 149972
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 154849 149834 154915 149837
rect 183502 149834 183508 149836
rect 154849 149832 183508 149834
rect 154849 149776 154854 149832
rect 154910 149776 183508 149832
rect 154849 149774 183508 149776
rect 154849 149771 154915 149774
rect 183502 149772 183508 149774
rect 183572 149772 183578 149836
rect 137277 149698 137343 149701
rect 142470 149698 142476 149700
rect 137277 149696 142476 149698
rect 137277 149640 137282 149696
rect 137338 149640 142476 149696
rect 137277 149638 142476 149640
rect 137277 149635 137343 149638
rect 142470 149636 142476 149638
rect 142540 149636 142546 149700
rect 151721 149698 151787 149701
rect 184974 149698 184980 149700
rect 151721 149696 184980 149698
rect 151721 149640 151726 149696
rect 151782 149640 184980 149696
rect 151721 149638 184980 149640
rect 151721 149635 151787 149638
rect 184974 149636 184980 149638
rect 185044 149636 185050 149700
rect 124949 148474 125015 148477
rect 145649 148474 145715 148477
rect 124949 148472 145715 148474
rect 124949 148416 124954 148472
rect 125010 148416 145654 148472
rect 145710 148416 145715 148472
rect 124949 148414 145715 148416
rect 124949 148411 125015 148414
rect 145649 148411 145715 148414
rect 100477 148338 100543 148341
rect 132677 148338 132743 148341
rect 100477 148336 132743 148338
rect 100477 148280 100482 148336
rect 100538 148280 132682 148336
rect 132738 148280 132743 148336
rect 100477 148278 132743 148280
rect 100477 148275 100543 148278
rect 132677 148275 132743 148278
rect 121913 147794 121979 147797
rect 122414 147794 122420 147796
rect 121913 147792 122420 147794
rect 121913 147736 121918 147792
rect 121974 147736 122420 147792
rect 121913 147734 122420 147736
rect 121913 147731 121979 147734
rect 122414 147732 122420 147734
rect 122484 147732 122490 147796
rect 201033 147794 201099 147797
rect 201166 147794 201172 147796
rect 201033 147792 201172 147794
rect 201033 147736 201038 147792
rect 201094 147736 201172 147792
rect 201033 147734 201172 147736
rect 201033 147731 201099 147734
rect 201166 147732 201172 147734
rect 201236 147732 201242 147796
rect 174169 147658 174235 147661
rect 193806 147658 193812 147660
rect 174169 147656 193812 147658
rect 174169 147600 174174 147656
rect 174230 147600 193812 147656
rect 174169 147598 193812 147600
rect 174169 147595 174235 147598
rect 193806 147596 193812 147598
rect 193876 147596 193882 147660
rect 174353 147522 174419 147525
rect 196382 147522 196388 147524
rect 174353 147520 196388 147522
rect 174353 147464 174358 147520
rect 174414 147464 196388 147520
rect 174353 147462 196388 147464
rect 174353 147459 174419 147462
rect 196382 147460 196388 147462
rect 196452 147460 196458 147524
rect 157425 147386 157491 147389
rect 181294 147386 181300 147388
rect 157425 147384 181300 147386
rect 157425 147328 157430 147384
rect 157486 147328 181300 147384
rect 157425 147326 181300 147328
rect 157425 147323 157491 147326
rect 181294 147324 181300 147326
rect 181364 147324 181370 147388
rect 172697 147250 172763 147253
rect 198038 147250 198044 147252
rect 172697 147248 198044 147250
rect 172697 147192 172702 147248
rect 172758 147192 198044 147248
rect 172697 147190 198044 147192
rect 172697 147187 172763 147190
rect 198038 147188 198044 147190
rect 198108 147188 198114 147252
rect 147581 147114 147647 147117
rect 180006 147114 180012 147116
rect 147581 147112 180012 147114
rect 147581 147056 147586 147112
rect 147642 147056 180012 147112
rect 147581 147054 180012 147056
rect 147581 147051 147647 147054
rect 180006 147052 180012 147054
rect 180076 147052 180082 147116
rect 117957 146978 118023 146981
rect 118417 146978 118483 146981
rect 117957 146976 118483 146978
rect 117957 146920 117962 146976
rect 118018 146920 118422 146976
rect 118478 146920 118483 146976
rect 117957 146918 118483 146920
rect 117957 146915 118023 146918
rect 118417 146915 118483 146918
rect 150617 146978 150683 146981
rect 183686 146978 183692 146980
rect 150617 146976 183692 146978
rect 150617 146920 150622 146976
rect 150678 146920 183692 146976
rect 150617 146918 183692 146920
rect 150617 146915 150683 146918
rect 183686 146916 183692 146918
rect 183756 146916 183762 146980
rect 195094 146916 195100 146980
rect 195164 146978 195170 146980
rect 195329 146978 195395 146981
rect 195164 146976 195395 146978
rect 195164 146920 195334 146976
rect 195390 146920 195395 146976
rect 195164 146918 195395 146920
rect 195164 146916 195170 146918
rect 195329 146915 195395 146918
rect 115422 146236 115428 146300
rect 115492 146298 115498 146300
rect 130285 146298 130351 146301
rect 115492 146296 130351 146298
rect 115492 146240 130290 146296
rect 130346 146240 130351 146296
rect 115492 146238 130351 146240
rect 115492 146236 115498 146238
rect 130285 146235 130351 146238
rect 197854 146236 197860 146300
rect 197924 146298 197930 146300
rect 198089 146298 198155 146301
rect 197924 146296 198155 146298
rect 197924 146240 198094 146296
rect 198150 146240 198155 146296
rect 197924 146238 198155 146240
rect 197924 146236 197930 146238
rect 198089 146235 198155 146238
rect 111558 146100 111564 146164
rect 111628 146162 111634 146164
rect 129825 146162 129891 146165
rect 111628 146160 129891 146162
rect 111628 146104 129830 146160
rect 129886 146104 129891 146160
rect 111628 146102 129891 146104
rect 111628 146100 111634 146102
rect 129825 146099 129891 146102
rect 174077 146162 174143 146165
rect 192518 146162 192524 146164
rect 174077 146160 192524 146162
rect 174077 146104 174082 146160
rect 174138 146104 192524 146160
rect 174077 146102 192524 146104
rect 174077 146099 174143 146102
rect 192518 146100 192524 146102
rect 192588 146100 192594 146164
rect 111190 145964 111196 146028
rect 111260 146026 111266 146028
rect 129733 146026 129799 146029
rect 111260 146024 129799 146026
rect 111260 145968 129738 146024
rect 129794 145968 129799 146024
rect 111260 145966 129799 145968
rect 111260 145964 111266 145966
rect 129733 145963 129799 145966
rect 175365 146026 175431 146029
rect 193990 146026 193996 146028
rect 175365 146024 193996 146026
rect 175365 145968 175370 146024
rect 175426 145968 193996 146024
rect 175365 145966 193996 145968
rect 175365 145963 175431 145966
rect 193990 145964 193996 145966
rect 194060 145964 194066 146028
rect 113766 145828 113772 145892
rect 113836 145890 113842 145892
rect 146661 145890 146727 145893
rect 113836 145888 146727 145890
rect 113836 145832 146666 145888
rect 146722 145832 146727 145888
rect 113836 145830 146727 145832
rect 113836 145828 113842 145830
rect 146661 145827 146727 145830
rect 175549 145890 175615 145893
rect 196566 145890 196572 145892
rect 175549 145888 196572 145890
rect 175549 145832 175554 145888
rect 175610 145832 196572 145888
rect 175549 145830 196572 145832
rect 175549 145827 175615 145830
rect 196566 145828 196572 145830
rect 196636 145828 196642 145892
rect 114134 145692 114140 145756
rect 114204 145754 114210 145756
rect 146293 145754 146359 145757
rect 114204 145752 146359 145754
rect 114204 145696 146298 145752
rect 146354 145696 146359 145752
rect 114204 145694 146359 145696
rect 114204 145692 114210 145694
rect 146293 145691 146359 145694
rect 158069 145754 158135 145757
rect 179822 145754 179828 145756
rect 158069 145752 179828 145754
rect 158069 145696 158074 145752
rect 158130 145696 179828 145752
rect 158069 145694 179828 145696
rect 158069 145691 158135 145694
rect 179822 145692 179828 145694
rect 179892 145692 179898 145756
rect 113950 145556 113956 145620
rect 114020 145618 114026 145620
rect 147673 145618 147739 145621
rect 114020 145616 147739 145618
rect 114020 145560 147678 145616
rect 147734 145560 147739 145616
rect 114020 145558 147739 145560
rect 114020 145556 114026 145558
rect 147673 145555 147739 145558
rect 164233 145618 164299 145621
rect 197670 145618 197676 145620
rect 164233 145616 197676 145618
rect 164233 145560 164238 145616
rect 164294 145560 197676 145616
rect 164233 145558 197676 145560
rect 164233 145555 164299 145558
rect 197670 145556 197676 145558
rect 197740 145556 197746 145620
rect 120758 144876 120764 144940
rect 120828 144938 120834 144940
rect 183829 144938 183895 144941
rect 120828 144936 183895 144938
rect 120828 144880 183834 144936
rect 183890 144880 183895 144936
rect 120828 144878 183895 144880
rect 120828 144876 120834 144878
rect 183829 144875 183895 144878
rect 193397 144938 193463 144941
rect 193622 144938 193628 144940
rect 193397 144936 193628 144938
rect 193397 144880 193402 144936
rect 193458 144880 193628 144936
rect 193397 144878 193628 144880
rect 193397 144875 193463 144878
rect 193622 144876 193628 144878
rect 193692 144876 193698 144940
rect 118182 144740 118188 144804
rect 118252 144802 118258 144804
rect 118325 144802 118391 144805
rect 118252 144800 118391 144802
rect 118252 144744 118330 144800
rect 118386 144744 118391 144800
rect 118252 144742 118391 144744
rect 118252 144740 118258 144742
rect 118325 144739 118391 144742
rect 168005 144802 168071 144805
rect 197486 144802 197492 144804
rect 168005 144800 197492 144802
rect 168005 144744 168010 144800
rect 168066 144744 197492 144800
rect 168005 144742 197492 144744
rect 168005 144739 168071 144742
rect 197486 144740 197492 144742
rect 197556 144740 197562 144804
rect 116301 144666 116367 144669
rect 144126 144666 144132 144668
rect 116301 144664 144132 144666
rect 116301 144608 116306 144664
rect 116362 144608 144132 144664
rect 116301 144606 144132 144608
rect 116301 144603 116367 144606
rect 144126 144604 144132 144606
rect 144196 144604 144202 144668
rect 166349 144666 166415 144669
rect 196198 144666 196204 144668
rect 166349 144664 196204 144666
rect 166349 144608 166354 144664
rect 166410 144608 196204 144664
rect 166349 144606 196204 144608
rect 166349 144603 166415 144606
rect 196198 144604 196204 144606
rect 196268 144604 196274 144668
rect 112662 144468 112668 144532
rect 112732 144530 112738 144532
rect 140865 144530 140931 144533
rect 112732 144528 140931 144530
rect 112732 144472 140870 144528
rect 140926 144472 140931 144528
rect 112732 144470 140931 144472
rect 112732 144468 112738 144470
rect 140865 144467 140931 144470
rect 162761 144530 162827 144533
rect 194542 144530 194548 144532
rect 162761 144528 194548 144530
rect 162761 144472 162766 144528
rect 162822 144472 194548 144528
rect 162761 144470 194548 144472
rect 162761 144467 162827 144470
rect 194542 144468 194548 144470
rect 194612 144468 194618 144532
rect 112846 144332 112852 144396
rect 112916 144394 112922 144396
rect 145833 144394 145899 144397
rect 112916 144392 145899 144394
rect 112916 144336 145838 144392
rect 145894 144336 145899 144392
rect 112916 144334 145899 144336
rect 112916 144332 112922 144334
rect 145833 144331 145899 144334
rect 160553 144394 160619 144397
rect 193438 144394 193444 144396
rect 160553 144392 193444 144394
rect 160553 144336 160558 144392
rect 160614 144336 193444 144392
rect 160553 144334 193444 144336
rect 160553 144331 160619 144334
rect 193438 144332 193444 144334
rect 193508 144332 193514 144396
rect 118182 144196 118188 144260
rect 118252 144258 118258 144260
rect 152549 144258 152615 144261
rect 118252 144256 152615 144258
rect 118252 144200 152554 144256
rect 152610 144200 152615 144256
rect 118252 144198 152615 144200
rect 118252 144196 118258 144198
rect 152549 144195 152615 144198
rect 156413 144258 156479 144261
rect 190494 144258 190500 144260
rect 156413 144256 190500 144258
rect 156413 144200 156418 144256
rect 156474 144200 190500 144256
rect 156413 144198 190500 144200
rect 156413 144195 156479 144198
rect 190494 144196 190500 144198
rect 190564 144196 190570 144260
rect 116710 144060 116716 144124
rect 116780 144122 116786 144124
rect 150985 144122 151051 144125
rect 116780 144120 151051 144122
rect 116780 144064 150990 144120
rect 151046 144064 151051 144120
rect 116780 144062 151051 144064
rect 116780 144060 116786 144062
rect 150985 144059 151051 144062
rect 158069 144122 158135 144125
rect 192150 144122 192156 144124
rect 158069 144120 192156 144122
rect 158069 144064 158074 144120
rect 158130 144064 192156 144120
rect 158069 144062 192156 144064
rect 158069 144059 158135 144062
rect 192150 144060 192156 144062
rect 192220 144060 192226 144124
rect 115606 143924 115612 143988
rect 115676 143986 115682 143988
rect 138657 143986 138723 143989
rect 115676 143984 138723 143986
rect 115676 143928 138662 143984
rect 138718 143928 138723 143984
rect 115676 143926 138723 143928
rect 115676 143924 115682 143926
rect 138657 143923 138723 143926
rect 163957 143986 164023 143989
rect 191966 143986 191972 143988
rect 163957 143984 191972 143986
rect 163957 143928 163962 143984
rect 164018 143928 191972 143984
rect 163957 143926 191972 143928
rect 163957 143923 164023 143926
rect 191966 143924 191972 143926
rect 192036 143924 192042 143988
rect 113030 143788 113036 143852
rect 113100 143850 113106 143852
rect 139393 143850 139459 143853
rect 113100 143848 139459 143850
rect 113100 143792 139398 143848
rect 139454 143792 139459 143848
rect 113100 143790 139459 143792
rect 113100 143788 113106 143790
rect 139393 143787 139459 143790
rect 165245 143442 165311 143445
rect 185945 143442 186011 143445
rect 187182 143442 187188 143444
rect 165245 143440 185226 143442
rect 165245 143384 165250 143440
rect 165306 143384 185226 143440
rect 165245 143382 185226 143384
rect 165245 143379 165311 143382
rect 111374 143244 111380 143308
rect 111444 143306 111450 143308
rect 132585 143306 132651 143309
rect 111444 143304 132651 143306
rect 111444 143248 132590 143304
rect 132646 143248 132651 143304
rect 111444 143246 132651 143248
rect 111444 143244 111450 143246
rect 132585 143243 132651 143246
rect 161933 143306 161999 143309
rect 185025 143306 185091 143309
rect 161933 143304 185091 143306
rect 161933 143248 161938 143304
rect 161994 143248 185030 143304
rect 185086 143248 185091 143304
rect 161933 143246 185091 143248
rect 185166 143306 185226 143382
rect 185945 143440 187188 143442
rect 185945 143384 185950 143440
rect 186006 143384 187188 143440
rect 185945 143382 187188 143384
rect 185945 143379 186011 143382
rect 187182 143380 187188 143382
rect 187252 143380 187258 143444
rect 189533 143306 189599 143309
rect 185166 143304 189599 143306
rect 185166 143248 189538 143304
rect 189594 143248 189599 143304
rect 185166 143246 189599 143248
rect 161933 143243 161999 143246
rect 185025 143243 185091 143246
rect 189533 143243 189599 143246
rect 121126 143108 121132 143172
rect 121196 143170 121202 143172
rect 145005 143170 145071 143173
rect 121196 143168 145071 143170
rect 121196 143112 145010 143168
rect 145066 143112 145071 143168
rect 121196 143110 145071 143112
rect 121196 143108 121202 143110
rect 145005 143107 145071 143110
rect 163589 143170 163655 143173
rect 191373 143170 191439 143173
rect 163589 143168 191439 143170
rect 163589 143112 163594 143168
rect 163650 143112 191378 143168
rect 191434 143112 191439 143168
rect 163589 143110 191439 143112
rect 163589 143107 163655 143110
rect 191373 143107 191439 143110
rect 121310 142972 121316 143036
rect 121380 143034 121386 143036
rect 148041 143034 148107 143037
rect 121380 143032 148107 143034
rect 121380 142976 148046 143032
rect 148102 142976 148107 143032
rect 121380 142974 148107 142976
rect 121380 142972 121386 142974
rect 148041 142971 148107 142974
rect 160001 143034 160067 143037
rect 190913 143034 190979 143037
rect 160001 143032 190979 143034
rect 160001 142976 160006 143032
rect 160062 142976 190918 143032
rect 190974 142976 190979 143032
rect 160001 142974 190979 142976
rect 160001 142971 160067 142974
rect 190913 142971 190979 142974
rect 119838 142836 119844 142900
rect 119908 142898 119914 142900
rect 146385 142898 146451 142901
rect 119908 142896 146451 142898
rect 119908 142840 146390 142896
rect 146446 142840 146451 142896
rect 119908 142838 146451 142840
rect 119908 142836 119914 142838
rect 146385 142835 146451 142838
rect 156965 142898 157031 142901
rect 189022 142898 189028 142900
rect 156965 142896 189028 142898
rect 156965 142840 156970 142896
rect 157026 142840 189028 142896
rect 156965 142838 189028 142840
rect 156965 142835 157031 142838
rect 189022 142836 189028 142838
rect 189092 142836 189098 142900
rect 119337 142762 119403 142765
rect 149697 142762 149763 142765
rect 119337 142760 149763 142762
rect 119337 142704 119342 142760
rect 119398 142704 149702 142760
rect 149758 142704 149763 142760
rect 119337 142702 149763 142704
rect 119337 142699 119403 142702
rect 149697 142699 149763 142702
rect 155309 142762 155375 142765
rect 185025 142762 185091 142765
rect 189574 142762 189580 142764
rect 155309 142760 180810 142762
rect 155309 142704 155314 142760
rect 155370 142704 180810 142760
rect 155309 142702 180810 142704
rect 155309 142699 155375 142702
rect 180750 142626 180810 142702
rect 185025 142760 189580 142762
rect 185025 142704 185030 142760
rect 185086 142704 189580 142760
rect 185025 142702 189580 142704
rect 185025 142699 185091 142702
rect 189574 142700 189580 142702
rect 189644 142700 189650 142764
rect 189206 142626 189212 142628
rect 180750 142566 189212 142626
rect 189206 142564 189212 142566
rect 189276 142564 189282 142628
rect 161381 142354 161447 142357
rect 161606 142354 161612 142356
rect 161336 142352 161612 142354
rect 161336 142296 161386 142352
rect 161442 142296 161612 142352
rect 161336 142294 161612 142296
rect 161381 142291 161447 142294
rect 161606 142292 161612 142294
rect 161676 142292 161682 142356
rect 120809 142218 120875 142221
rect 122966 142218 122972 142220
rect 120809 142216 122972 142218
rect 120809 142160 120814 142216
rect 120870 142160 122972 142216
rect 120809 142158 122972 142160
rect 120809 142155 120875 142158
rect 122966 142156 122972 142158
rect 123036 142218 123042 142220
rect 124029 142218 124095 142221
rect 123036 142216 124095 142218
rect 123036 142160 124034 142216
rect 124090 142160 124095 142216
rect 123036 142158 124095 142160
rect 123036 142156 123042 142158
rect 124029 142155 124095 142158
rect 153653 142218 153719 142221
rect 178217 142218 178283 142221
rect 153653 142216 178283 142218
rect 153653 142160 153658 142216
rect 153714 142160 178222 142216
rect 178278 142160 178283 142216
rect 153653 142158 178283 142160
rect 153653 142155 153719 142158
rect 178217 142155 178283 142158
rect 161473 142082 161539 142085
rect 191782 142082 191788 142084
rect 161473 142080 191788 142082
rect 161473 142024 161478 142080
rect 161534 142024 191788 142080
rect 161473 142022 191788 142024
rect 161473 142019 161539 142022
rect 191782 142020 191788 142022
rect 191852 142020 191858 142084
rect 117078 141748 117084 141812
rect 117148 141810 117154 141812
rect 140313 141810 140379 141813
rect 117148 141808 140379 141810
rect 117148 141752 140318 141808
rect 140374 141752 140379 141808
rect 117148 141750 140379 141752
rect 117148 141748 117154 141750
rect 140313 141747 140379 141750
rect 118366 141612 118372 141676
rect 118436 141674 118442 141676
rect 142245 141674 142311 141677
rect 118436 141672 142311 141674
rect 118436 141616 142250 141672
rect 142306 141616 142311 141672
rect 118436 141614 142311 141616
rect 118436 141612 118442 141614
rect 142245 141611 142311 141614
rect 116894 141476 116900 141540
rect 116964 141538 116970 141540
rect 143625 141538 143691 141541
rect 116964 141536 143691 141538
rect 116964 141480 143630 141536
rect 143686 141480 143691 141536
rect 116964 141478 143691 141480
rect 116964 141476 116970 141478
rect 143625 141475 143691 141478
rect 180149 141538 180215 141541
rect 190494 141538 190500 141540
rect 180149 141536 190500 141538
rect 180149 141480 180154 141536
rect 180210 141480 190500 141536
rect 180149 141478 190500 141480
rect 180149 141475 180215 141478
rect 190494 141476 190500 141478
rect 190564 141476 190570 141540
rect 115790 141340 115796 141404
rect 115860 141402 115866 141404
rect 150433 141402 150499 141405
rect 115860 141400 150499 141402
rect 115860 141344 150438 141400
rect 150494 141344 150499 141400
rect 115860 141342 150499 141344
rect 115860 141340 115866 141342
rect 150433 141339 150499 141342
rect 162853 141402 162919 141405
rect 183870 141402 183876 141404
rect 162853 141400 183876 141402
rect 162853 141344 162858 141400
rect 162914 141344 183876 141400
rect 162853 141342 183876 141344
rect 162853 141339 162919 141342
rect 183870 141340 183876 141342
rect 183940 141340 183946 141404
rect 141366 141204 141372 141268
rect 141436 141266 141442 141268
rect 141509 141266 141575 141269
rect 141436 141264 141575 141266
rect 141436 141208 141514 141264
rect 141570 141208 141575 141264
rect 141436 141206 141575 141208
rect 141436 141204 141442 141206
rect 141509 141203 141575 141206
rect 176653 141266 176719 141269
rect 177798 141266 177804 141268
rect 176653 141264 177804 141266
rect 176653 141208 176658 141264
rect 176714 141208 177804 141264
rect 176653 141206 177804 141208
rect 176653 141203 176719 141206
rect 177798 141204 177804 141206
rect 177868 141204 177874 141268
rect 141417 141130 141483 141133
rect 141550 141130 141556 141132
rect 141417 141128 141556 141130
rect 141417 141072 141422 141128
rect 141478 141072 141556 141128
rect 141417 141070 141556 141072
rect 141417 141067 141483 141070
rect 141550 141068 141556 141070
rect 141620 141068 141626 141132
rect 176745 141130 176811 141133
rect 177430 141130 177436 141132
rect 176745 141128 177436 141130
rect 176745 141072 176750 141128
rect 176806 141072 177436 141128
rect 176745 141070 177436 141072
rect 176745 141067 176811 141070
rect 177430 141068 177436 141070
rect 177500 141068 177506 141132
rect 126237 140994 126303 140997
rect 188286 140994 188292 140996
rect 126237 140992 188292 140994
rect 126237 140936 126242 140992
rect 126298 140936 188292 140992
rect 126237 140934 188292 140936
rect 126237 140931 126303 140934
rect 188286 140932 188292 140934
rect 188356 140932 188362 140996
rect 125501 140858 125567 140861
rect 192334 140858 192340 140860
rect 125501 140856 192340 140858
rect 125501 140800 125506 140856
rect 125562 140800 192340 140856
rect 125501 140798 192340 140800
rect 125501 140795 125567 140798
rect 192334 140796 192340 140798
rect 192404 140796 192410 140860
rect 180793 140722 180859 140725
rect 181161 140722 181227 140725
rect 183921 140722 183987 140725
rect 184749 140722 184815 140725
rect 190821 140724 190887 140725
rect 190821 140722 190868 140724
rect 180793 140720 181227 140722
rect 180793 140664 180798 140720
rect 180854 140664 181166 140720
rect 181222 140664 181227 140720
rect 180793 140662 181227 140664
rect 180793 140659 180859 140662
rect 181161 140659 181227 140662
rect 183142 140720 184815 140722
rect 183142 140664 183926 140720
rect 183982 140664 184754 140720
rect 184810 140664 184815 140720
rect 183142 140662 184815 140664
rect 190776 140720 190868 140722
rect 190776 140664 190826 140720
rect 190776 140662 190868 140664
rect 120574 140524 120580 140588
rect 120644 140586 120650 140588
rect 183142 140586 183202 140662
rect 183921 140659 183987 140662
rect 184749 140659 184815 140662
rect 190821 140660 190868 140662
rect 190932 140660 190938 140724
rect 190821 140659 190887 140660
rect 185853 140586 185919 140589
rect 120644 140526 183202 140586
rect 184062 140584 185919 140586
rect 184062 140528 185858 140584
rect 185914 140528 185919 140584
rect 184062 140526 185919 140528
rect 120644 140524 120650 140526
rect 116526 140388 116532 140452
rect 116596 140450 116602 140452
rect 184062 140450 184122 140526
rect 185853 140523 185919 140526
rect 184381 140452 184447 140453
rect 184381 140450 184428 140452
rect 116596 140390 184122 140450
rect 184336 140448 184428 140450
rect 184336 140392 184386 140448
rect 184336 140390 184428 140392
rect 116596 140388 116602 140390
rect 184381 140388 184428 140390
rect 184492 140388 184498 140452
rect 184381 140387 184447 140388
rect 123477 140314 123543 140317
rect 126605 140314 126671 140317
rect 123477 140312 126671 140314
rect 123477 140256 123482 140312
rect 123538 140256 126610 140312
rect 126666 140256 126671 140312
rect 123477 140254 126671 140256
rect 123477 140251 123543 140254
rect 126605 140251 126671 140254
rect 170029 140314 170095 140317
rect 191598 140314 191604 140316
rect 170029 140312 191604 140314
rect 170029 140256 170034 140312
rect 170090 140256 191604 140312
rect 170029 140254 191604 140256
rect 170029 140251 170095 140254
rect 191598 140252 191604 140254
rect 191668 140252 191674 140316
rect 122230 140116 122236 140180
rect 122300 140178 122306 140180
rect 127617 140178 127683 140181
rect 122300 140176 127683 140178
rect 122300 140120 127622 140176
rect 127678 140120 127683 140176
rect 122300 140118 127683 140120
rect 122300 140116 122306 140118
rect 127617 140115 127683 140118
rect 156505 140178 156571 140181
rect 171225 140178 171291 140181
rect 156505 140176 171291 140178
rect 156505 140120 156510 140176
rect 156566 140120 171230 140176
rect 171286 140120 171291 140176
rect 156505 140118 171291 140120
rect 156505 140115 156571 140118
rect 171225 140115 171291 140118
rect 178033 140178 178099 140181
rect 188470 140178 188476 140180
rect 178033 140176 188476 140178
rect 178033 140120 178038 140176
rect 178094 140120 188476 140176
rect 178033 140118 188476 140120
rect 178033 140115 178099 140118
rect 188470 140116 188476 140118
rect 188540 140116 188546 140180
rect 154757 140042 154823 140045
rect 178902 140042 178908 140044
rect 154757 140040 178908 140042
rect 154757 139984 154762 140040
rect 154818 139984 178908 140040
rect 154757 139982 178908 139984
rect 154757 139979 154823 139982
rect 178902 139980 178908 139982
rect 178972 139980 178978 140044
rect 179137 140042 179203 140045
rect 179137 140040 190470 140042
rect 179137 139984 179142 140040
rect 179198 139984 190470 140040
rect 179137 139982 190470 139984
rect 179137 139979 179203 139982
rect 119286 139844 119292 139908
rect 119356 139906 119362 139908
rect 181805 139906 181871 139909
rect 189574 139906 189580 139908
rect 119356 139846 180810 139906
rect 119356 139844 119362 139846
rect 171225 139770 171291 139773
rect 178534 139770 178540 139772
rect 171225 139768 178540 139770
rect 171225 139712 171230 139768
rect 171286 139712 178540 139768
rect 171225 139710 178540 139712
rect 171225 139707 171291 139710
rect 178534 139708 178540 139710
rect 178604 139708 178610 139772
rect 180750 139770 180810 139846
rect 181805 139904 189580 139906
rect 181805 139848 181810 139904
rect 181866 139848 189580 139904
rect 181805 139846 189580 139848
rect 181805 139843 181871 139846
rect 189574 139844 189580 139846
rect 189644 139844 189650 139908
rect 190410 139906 190470 139982
rect 191966 139906 191972 139908
rect 190410 139846 191972 139906
rect 191966 139844 191972 139846
rect 192036 139844 192042 139908
rect 181897 139770 181963 139773
rect 185761 139772 185827 139773
rect 180750 139768 181963 139770
rect 180750 139712 181902 139768
rect 181958 139712 181963 139768
rect 180750 139710 181963 139712
rect 181897 139707 181963 139710
rect 185710 139708 185716 139772
rect 185780 139770 185827 139772
rect 185780 139768 185872 139770
rect 185822 139712 185872 139768
rect 185780 139710 185872 139712
rect 185780 139708 185827 139710
rect 189022 139708 189028 139772
rect 189092 139770 189098 139772
rect 189809 139770 189875 139773
rect 189092 139768 189875 139770
rect 189092 139712 189814 139768
rect 189870 139712 189875 139768
rect 189092 139710 189875 139712
rect 189092 139708 189098 139710
rect 185761 139707 185827 139708
rect 189809 139707 189875 139710
rect 123201 139634 123267 139637
rect 125041 139634 125107 139637
rect 123201 139632 125107 139634
rect 123201 139576 123206 139632
rect 123262 139576 125046 139632
rect 125102 139576 125107 139632
rect 123201 139574 125107 139576
rect 123201 139571 123267 139574
rect 125041 139571 125107 139574
rect 181897 139634 181963 139637
rect 289077 139634 289143 139637
rect 181897 139632 289143 139634
rect 181897 139576 181902 139632
rect 181958 139576 289082 139632
rect 289138 139576 289143 139632
rect 181897 139574 289143 139576
rect 181897 139571 181963 139574
rect 289077 139571 289143 139574
rect 31017 139498 31083 139501
rect 181253 139498 181319 139501
rect 31017 139496 181319 139498
rect 31017 139440 31022 139496
rect 31078 139440 181258 139496
rect 181314 139440 181319 139496
rect 31017 139438 181319 139440
rect 31017 139435 31083 139438
rect 181253 139435 181319 139438
rect 182817 139498 182883 139501
rect 183318 139498 183324 139500
rect 182817 139496 183324 139498
rect 182817 139440 182822 139496
rect 182878 139440 183324 139496
rect 182817 139438 183324 139440
rect 182817 139435 182883 139438
rect 183318 139436 183324 139438
rect 183388 139436 183394 139500
rect 184657 139498 184723 139501
rect 576117 139498 576183 139501
rect 184657 139496 576183 139498
rect 184657 139440 184662 139496
rect 184718 139440 576122 139496
rect 576178 139440 576183 139496
rect 184657 139438 576183 139440
rect 184657 139435 184723 139438
rect 576117 139435 576183 139438
rect 122046 139300 122052 139364
rect 122116 139362 122122 139364
rect 124949 139362 125015 139365
rect 126145 139362 126211 139365
rect 122116 139360 125015 139362
rect 122116 139304 124954 139360
rect 125010 139304 125015 139360
rect 122116 139302 125015 139304
rect 122116 139300 122122 139302
rect 124949 139299 125015 139302
rect 125182 139360 126211 139362
rect 125182 139304 126150 139360
rect 126206 139304 126211 139360
rect 125182 139302 126211 139304
rect 115105 139090 115171 139093
rect 125182 139090 125242 139302
rect 126145 139299 126211 139302
rect 126278 139300 126284 139364
rect 126348 139362 126354 139364
rect 126697 139362 126763 139365
rect 126348 139360 126763 139362
rect 126348 139304 126702 139360
rect 126758 139304 126763 139360
rect 126348 139302 126763 139304
rect 126348 139300 126354 139302
rect 126697 139299 126763 139302
rect 127934 139300 127940 139364
rect 128004 139362 128010 139364
rect 128261 139362 128327 139365
rect 128004 139360 128327 139362
rect 128004 139304 128266 139360
rect 128322 139304 128327 139360
rect 128004 139302 128327 139304
rect 128004 139300 128010 139302
rect 128261 139299 128327 139302
rect 131982 139300 131988 139364
rect 132052 139362 132058 139364
rect 132217 139362 132283 139365
rect 133045 139362 133111 139365
rect 145741 139362 145807 139365
rect 132052 139360 132283 139362
rect 132052 139304 132222 139360
rect 132278 139304 132283 139360
rect 132052 139302 132283 139304
rect 132052 139300 132058 139302
rect 132217 139299 132283 139302
rect 132450 139360 133111 139362
rect 132450 139304 133050 139360
rect 133106 139304 133111 139360
rect 132450 139302 133111 139304
rect 115105 139088 125242 139090
rect 115105 139032 115110 139088
rect 115166 139032 125242 139088
rect 115105 139030 125242 139032
rect 115105 139027 115171 139030
rect 113725 138954 113791 138957
rect 132450 138954 132510 139302
rect 133045 139299 133111 139302
rect 142110 139360 145807 139362
rect 142110 139304 145746 139360
rect 145802 139304 145807 139360
rect 142110 139302 145807 139304
rect 113725 138952 132510 138954
rect 113725 138896 113730 138952
rect 113786 138896 132510 138952
rect 113725 138894 132510 138896
rect 113725 138891 113791 138894
rect 123293 138818 123359 138821
rect 142110 138818 142170 139302
rect 145741 139299 145807 139302
rect 150750 139300 150756 139364
rect 150820 139362 150826 139364
rect 150893 139362 150959 139365
rect 154021 139362 154087 139365
rect 150820 139360 150959 139362
rect 150820 139304 150898 139360
rect 150954 139304 150959 139360
rect 150820 139302 150959 139304
rect 150820 139300 150826 139302
rect 150893 139299 150959 139302
rect 151770 139360 154087 139362
rect 151770 139304 154026 139360
rect 154082 139304 154087 139360
rect 151770 139302 154087 139304
rect 123293 138816 142170 138818
rect 123293 138760 123298 138816
rect 123354 138760 142170 138816
rect 123293 138758 142170 138760
rect 123293 138755 123359 138758
rect 119613 138682 119679 138685
rect 151770 138682 151830 139302
rect 154021 139299 154087 139302
rect 155350 139300 155356 139364
rect 155420 139362 155426 139364
rect 155677 139362 155743 139365
rect 155420 139360 155743 139362
rect 155420 139304 155682 139360
rect 155738 139304 155743 139360
rect 155420 139302 155743 139304
rect 155420 139300 155426 139302
rect 155677 139299 155743 139302
rect 155861 139362 155927 139365
rect 157057 139362 157123 139365
rect 155861 139360 155970 139362
rect 155861 139304 155866 139360
rect 155922 139304 155970 139360
rect 155861 139299 155970 139304
rect 157057 139360 157258 139362
rect 157057 139304 157062 139360
rect 157118 139304 157258 139360
rect 157057 139302 157258 139304
rect 157057 139299 157123 139302
rect 154798 139164 154804 139228
rect 154868 139226 154874 139228
rect 155910 139226 155970 139299
rect 154868 139166 155970 139226
rect 157198 139226 157258 139302
rect 159214 139300 159220 139364
rect 159284 139362 159290 139364
rect 159541 139362 159607 139365
rect 159284 139360 159607 139362
rect 159284 139304 159546 139360
rect 159602 139304 159607 139360
rect 159284 139302 159607 139304
rect 159284 139300 159290 139302
rect 159541 139299 159607 139302
rect 159725 139362 159791 139365
rect 159950 139362 159956 139364
rect 159725 139360 159956 139362
rect 159725 139304 159730 139360
rect 159786 139304 159956 139360
rect 159725 139302 159956 139304
rect 159725 139299 159791 139302
rect 159950 139300 159956 139302
rect 160020 139300 160026 139364
rect 178401 139360 178467 139365
rect 178401 139304 178406 139360
rect 178462 139304 178467 139360
rect 178401 139299 178467 139304
rect 178861 139362 178927 139365
rect 180241 139362 180307 139365
rect 188245 139362 188311 139365
rect 178861 139360 178970 139362
rect 178861 139304 178866 139360
rect 178922 139304 178970 139360
rect 178861 139299 178970 139304
rect 180241 139360 188311 139362
rect 180241 139304 180246 139360
rect 180302 139304 188250 139360
rect 188306 139304 188311 139360
rect 180241 139302 188311 139304
rect 180241 139299 180307 139302
rect 188245 139299 188311 139302
rect 580441 139362 580507 139365
rect 583520 139362 584960 139452
rect 580441 139360 584960 139362
rect 580441 139304 580446 139360
rect 580502 139304 584960 139360
rect 580441 139302 584960 139304
rect 580441 139299 580507 139302
rect 157198 139166 161490 139226
rect 154868 139164 154874 139166
rect 119613 138680 151830 138682
rect 119613 138624 119618 138680
rect 119674 138624 151830 138680
rect 119613 138622 151830 138624
rect 161430 138682 161490 139166
rect 178404 138818 178464 139299
rect 178910 139226 178970 139299
rect 187325 139226 187391 139229
rect 178910 139224 187391 139226
rect 178910 139168 187330 139224
rect 187386 139168 187391 139224
rect 583520 139212 584960 139302
rect 178910 139166 187391 139168
rect 187325 139163 187391 139166
rect 185710 139028 185716 139092
rect 185780 139090 185786 139092
rect 194961 139090 195027 139093
rect 185780 139088 195027 139090
rect 185780 139032 194966 139088
rect 195022 139032 195027 139088
rect 185780 139030 195027 139032
rect 185780 139028 185786 139030
rect 194961 139027 195027 139030
rect 183318 138892 183324 138956
rect 183388 138954 183394 138956
rect 193397 138954 193463 138957
rect 183388 138952 193463 138954
rect 183388 138896 193402 138952
rect 193458 138896 193463 138952
rect 183388 138894 193463 138896
rect 183388 138892 183394 138894
rect 193397 138891 193463 138894
rect 178404 138758 190470 138818
rect 190410 138682 190470 138758
rect 190821 138682 190887 138685
rect 161430 138622 180810 138682
rect 190410 138680 190887 138682
rect 190410 138624 190826 138680
rect 190882 138624 190887 138680
rect 190410 138622 190887 138624
rect 119613 138619 119679 138622
rect 180750 138546 180810 138622
rect 190821 138619 190887 138622
rect 191097 138546 191163 138549
rect 180750 138544 191163 138546
rect 180750 138488 191102 138544
rect 191158 138488 191163 138544
rect 180750 138486 191163 138488
rect 191097 138483 191163 138486
rect 184422 138348 184428 138412
rect 184492 138410 184498 138412
rect 192293 138410 192359 138413
rect 184492 138408 192359 138410
rect 184492 138352 192298 138408
rect 192354 138352 192359 138408
rect 184492 138350 192359 138352
rect 184492 138348 184498 138350
rect 192293 138347 192359 138350
rect 186262 138212 186268 138276
rect 186332 138274 186338 138276
rect 187509 138274 187575 138277
rect 186332 138272 187575 138274
rect 186332 138216 187514 138272
rect 187570 138216 187575 138272
rect 186332 138214 187575 138216
rect 186332 138212 186338 138214
rect 187509 138211 187575 138214
rect 187182 138076 187188 138140
rect 187252 138138 187258 138140
rect 187417 138138 187483 138141
rect 187252 138136 187483 138138
rect 187252 138080 187422 138136
rect 187478 138080 187483 138136
rect 187252 138078 187483 138080
rect 187252 138076 187258 138078
rect 187417 138075 187483 138078
rect 122230 137940 122236 138004
rect 122300 138002 122306 138004
rect 122782 138002 122788 138004
rect 122300 137942 122788 138002
rect 122300 137940 122306 137942
rect 122782 137940 122788 137942
rect 122852 137940 122858 138004
rect 185342 137940 185348 138004
rect 185412 138002 185418 138004
rect 196525 138002 196591 138005
rect 185412 138000 196591 138002
rect 185412 137944 196530 138000
rect 196586 137944 196591 138000
rect 185412 137942 196591 137944
rect 185412 137940 185418 137942
rect 196525 137939 196591 137942
rect 185158 137804 185164 137868
rect 185228 137866 185234 137868
rect 198089 137866 198155 137869
rect 185228 137864 198155 137866
rect 185228 137808 198094 137864
rect 198150 137808 198155 137864
rect 185228 137806 198155 137808
rect 185228 137804 185234 137806
rect 198089 137803 198155 137806
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 122189 128482 122255 128485
rect 122782 128482 122788 128484
rect 122189 128480 122788 128482
rect 122189 128424 122194 128480
rect 122250 128424 122788 128480
rect 122189 128422 122788 128424
rect 122189 128419 122255 128422
rect 122782 128420 122788 128422
rect 122852 128420 122858 128484
rect 186078 127604 186084 127668
rect 186148 127666 186154 127668
rect 188521 127666 188587 127669
rect 186148 127664 188587 127666
rect 186148 127608 188526 127664
rect 188582 127608 188587 127664
rect 186148 127606 188587 127608
rect 186148 127604 186154 127606
rect 188521 127603 188587 127606
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 188470 125564 188476 125628
rect 188540 125626 188546 125628
rect 583526 125626 583586 125838
rect 188540 125566 583586 125626
rect 188540 125564 188546 125566
rect -960 123572 480 123812
rect 122189 123178 122255 123181
rect 122782 123178 122788 123180
rect 122189 123176 122788 123178
rect 122189 123120 122194 123176
rect 122250 123120 122788 123176
rect 122189 123118 122788 123120
rect 122189 123115 122255 123118
rect 122782 123116 122788 123118
rect 122852 123116 122858 123180
rect 121913 122770 121979 122773
rect 122097 122770 122163 122773
rect 121913 122768 122163 122770
rect 121913 122712 121918 122768
rect 121974 122712 122102 122768
rect 122158 122712 122163 122768
rect 121913 122710 122163 122712
rect 121913 122707 121979 122710
rect 122097 122707 122163 122710
rect 122189 122498 122255 122501
rect 122782 122498 122788 122500
rect 122189 122496 122788 122498
rect 122189 122440 122194 122496
rect 122250 122440 122788 122496
rect 122189 122438 122788 122440
rect 122189 122435 122255 122438
rect 122782 122436 122788 122438
rect 122852 122436 122858 122500
rect 122189 113522 122255 113525
rect 122782 113522 122788 113524
rect 122189 113520 122788 113522
rect 122189 113464 122194 113520
rect 122250 113464 122788 113520
rect 122189 113462 122788 113464
rect 122189 113459 122255 113462
rect 122782 113460 122788 113462
rect 122852 113460 122858 113524
rect 121913 113386 121979 113389
rect 121913 113384 122114 113386
rect 121913 113328 121918 113384
rect 121974 113328 122114 113384
rect 121913 113326 122114 113328
rect 121913 113323 121979 113326
rect 122054 113253 122114 113326
rect 122054 113248 122163 113253
rect 122054 113192 122102 113248
rect 122158 113192 122163 113248
rect 122054 113190 122163 113192
rect 122097 113187 122163 113190
rect 122189 112842 122255 112845
rect 122782 112842 122788 112844
rect 122189 112840 122788 112842
rect 122189 112784 122194 112840
rect 122250 112784 122788 112840
rect 122189 112782 122788 112784
rect 122189 112779 122255 112782
rect 122782 112780 122788 112782
rect 122852 112780 122858 112844
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 189574 111828 189580 111892
rect 189644 111890 189650 111892
rect 583526 111890 583586 112646
rect 189644 111830 583586 111890
rect 189644 111828 189650 111830
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 122189 103866 122255 103869
rect 122782 103866 122788 103868
rect 122189 103864 122788 103866
rect 122189 103808 122194 103864
rect 122250 103808 122788 103864
rect 122189 103806 122788 103808
rect 122189 103803 122255 103806
rect 122782 103804 122788 103806
rect 122852 103804 122858 103868
rect 122097 103458 122163 103461
rect 122054 103456 122163 103458
rect 122054 103400 122102 103456
rect 122158 103400 122163 103456
rect 122054 103395 122163 103400
rect 121913 103322 121979 103325
rect 122054 103322 122114 103395
rect 121913 103320 122114 103322
rect 121913 103264 121918 103320
rect 121974 103264 122114 103320
rect 121913 103262 122114 103264
rect 121913 103259 121979 103262
rect 122189 103186 122255 103189
rect 122782 103186 122788 103188
rect 122189 103184 122788 103186
rect 122189 103128 122194 103184
rect 122250 103128 122788 103184
rect 122189 103126 122788 103128
rect 122189 103123 122255 103126
rect 122782 103124 122788 103126
rect 122852 103124 122858 103188
rect 580257 99514 580323 99517
rect 583520 99514 584960 99604
rect 580257 99512 584960 99514
rect 580257 99456 580262 99512
rect 580318 99456 584960 99512
rect 580257 99454 584960 99456
rect 580257 99451 580323 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 122189 94210 122255 94213
rect 122782 94210 122788 94212
rect 122189 94208 122788 94210
rect 122189 94152 122194 94208
rect 122250 94152 122788 94208
rect 122189 94150 122788 94152
rect 122189 94147 122255 94150
rect 122782 94148 122788 94150
rect 122852 94148 122858 94212
rect 121913 94074 121979 94077
rect 121913 94072 122114 94074
rect 121913 94016 121918 94072
rect 121974 94016 122114 94072
rect 121913 94014 122114 94016
rect 121913 94011 121979 94014
rect 122054 93941 122114 94014
rect 122054 93936 122163 93941
rect 122054 93880 122102 93936
rect 122158 93880 122163 93936
rect 122054 93878 122163 93880
rect 122097 93875 122163 93878
rect 122189 93530 122255 93533
rect 122782 93530 122788 93532
rect 122189 93528 122788 93530
rect 122189 93472 122194 93528
rect 122250 93472 122788 93528
rect 122189 93470 122788 93472
rect 122189 93467 122255 93470
rect 122782 93468 122788 93470
rect 122852 93468 122858 93532
rect 122189 89722 122255 89725
rect 122782 89722 122788 89724
rect 122189 89720 122788 89722
rect 122189 89664 122194 89720
rect 122250 89664 122788 89720
rect 122189 89662 122788 89664
rect 122189 89659 122255 89662
rect 122782 89660 122788 89662
rect 122852 89660 122858 89724
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 121637 85234 121703 85237
rect 122005 85234 122071 85237
rect 121637 85232 122071 85234
rect 121637 85176 121642 85232
rect 121698 85176 122010 85232
rect 122066 85176 122071 85232
rect 121637 85174 122071 85176
rect 121637 85171 121703 85174
rect 122005 85171 122071 85174
rect 122373 85098 122439 85101
rect 122373 85096 122482 85098
rect 122373 85040 122378 85096
rect 122434 85040 122482 85096
rect 122373 85035 122482 85040
rect -960 84690 480 84780
rect 122422 84693 122482 85035
rect -960 84630 6930 84690
rect -960 84540 480 84630
rect 6870 84282 6930 84630
rect 122373 84688 122482 84693
rect 122373 84632 122378 84688
rect 122434 84632 122482 84688
rect 122373 84630 122482 84632
rect 122373 84627 122439 84630
rect 119286 84282 119292 84284
rect 6870 84222 119292 84282
rect 119286 84220 119292 84222
rect 119356 84220 119362 84284
rect 134558 81908 134564 81972
rect 134628 81970 134634 81972
rect 135110 81970 135116 81972
rect 134628 81910 135116 81970
rect 134628 81908 134634 81910
rect 135110 81908 135116 81910
rect 135180 81908 135186 81972
rect 95233 81562 95299 81565
rect 139342 81562 139348 81564
rect 95233 81560 139348 81562
rect 95233 81504 95238 81560
rect 95294 81504 139348 81560
rect 95233 81502 139348 81504
rect 95233 81499 95299 81502
rect 139342 81500 139348 81502
rect 139412 81500 139418 81564
rect 137318 81364 137324 81428
rect 137388 81426 137394 81428
rect 142838 81426 142844 81428
rect 137388 81366 142844 81426
rect 137388 81364 137394 81366
rect 142838 81364 142844 81366
rect 142908 81364 142914 81428
rect 130694 81228 130700 81292
rect 130764 81290 130770 81292
rect 143206 81290 143212 81292
rect 130764 81230 143212 81290
rect 130764 81228 130770 81230
rect 143206 81228 143212 81230
rect 143276 81228 143282 81292
rect 176510 81228 176516 81292
rect 176580 81290 176586 81292
rect 195329 81290 195395 81293
rect 176580 81288 195395 81290
rect 176580 81232 195334 81288
rect 195390 81232 195395 81288
rect 176580 81230 195395 81232
rect 176580 81228 176586 81230
rect 195329 81227 195395 81230
rect 130510 81092 130516 81156
rect 130580 81154 130586 81156
rect 143390 81154 143396 81156
rect 130580 81094 143396 81154
rect 130580 81092 130586 81094
rect 143390 81092 143396 81094
rect 143460 81092 143466 81156
rect 173198 81092 173204 81156
rect 173268 81154 173274 81156
rect 195513 81154 195579 81157
rect 173268 81152 195579 81154
rect 173268 81096 195518 81152
rect 195574 81096 195579 81152
rect 173268 81094 195579 81096
rect 173268 81092 173274 81094
rect 195513 81091 195579 81094
rect 127934 80956 127940 81020
rect 128004 81018 128010 81020
rect 147990 81018 147996 81020
rect 128004 80958 147996 81018
rect 128004 80956 128010 80958
rect 147990 80956 147996 80958
rect 148060 80956 148066 81020
rect 175222 80956 175228 81020
rect 175292 81018 175298 81020
rect 197077 81018 197143 81021
rect 175292 81016 197143 81018
rect 175292 80960 197082 81016
rect 197138 80960 197143 81016
rect 175292 80958 197143 80960
rect 175292 80956 175298 80958
rect 197077 80955 197143 80958
rect 124990 80820 124996 80884
rect 125060 80882 125066 80884
rect 144862 80882 144868 80884
rect 125060 80822 144868 80882
rect 125060 80820 125066 80822
rect 144862 80820 144868 80822
rect 144932 80820 144938 80884
rect 160318 80820 160324 80884
rect 160388 80882 160394 80884
rect 199101 80882 199167 80885
rect 523125 80882 523191 80885
rect 160388 80822 177636 80882
rect 160388 80820 160394 80822
rect 116393 80746 116459 80749
rect 116393 80744 138030 80746
rect 116393 80688 116398 80744
rect 116454 80688 138030 80744
rect 116393 80686 138030 80688
rect 116393 80683 116459 80686
rect 131941 80610 132007 80613
rect 132166 80610 132172 80612
rect 131941 80608 132172 80610
rect 131941 80552 131946 80608
rect 132002 80552 132172 80608
rect 131941 80550 132172 80552
rect 131941 80547 132007 80550
rect 132166 80548 132172 80550
rect 132236 80548 132242 80612
rect 137970 80610 138030 80686
rect 170438 80684 170444 80748
rect 170508 80746 170514 80748
rect 170508 80686 172530 80746
rect 170508 80684 170514 80686
rect 137970 80550 147874 80610
rect 145046 80474 145052 80476
rect 137970 80414 145052 80474
rect 122465 80338 122531 80341
rect 122782 80338 122788 80340
rect 122465 80336 122788 80338
rect 122465 80280 122470 80336
rect 122526 80280 122788 80336
rect 122465 80278 122788 80280
rect 122465 80275 122531 80278
rect 122782 80276 122788 80278
rect 122852 80276 122858 80340
rect 126278 80276 126284 80340
rect 126348 80338 126354 80340
rect 130929 80338 130995 80341
rect 137970 80338 138030 80414
rect 145046 80412 145052 80414
rect 145116 80412 145122 80476
rect 126348 80336 138030 80338
rect 126348 80280 130934 80336
rect 130990 80280 138030 80336
rect 126348 80278 138030 80280
rect 126348 80276 126354 80278
rect 130929 80275 130995 80278
rect 138238 80276 138244 80340
rect 138308 80338 138314 80340
rect 138308 80278 146356 80338
rect 138308 80276 138314 80278
rect 105721 80202 105787 80205
rect 105721 80200 139410 80202
rect 105721 80144 105726 80200
rect 105782 80144 139410 80200
rect 105721 80142 139410 80144
rect 105721 80139 105787 80142
rect 122966 80004 122972 80068
rect 123036 80066 123042 80068
rect 131849 80066 131915 80069
rect 123036 80064 131915 80066
rect 123036 80008 131854 80064
rect 131910 80008 131915 80064
rect 123036 80006 131915 80008
rect 123036 80004 123042 80006
rect 131849 80003 131915 80006
rect 134374 80004 134380 80068
rect 134444 80066 134450 80068
rect 134444 80006 134902 80066
rect 134444 80004 134450 80006
rect 132539 79962 132605 79967
rect 132999 79964 133065 79967
rect 130193 79930 130259 79933
rect 132539 79930 132544 79962
rect 130193 79928 132544 79930
rect 130193 79872 130198 79928
rect 130254 79906 132544 79928
rect 132600 79906 132605 79962
rect 132956 79962 133065 79964
rect 130254 79901 132605 79906
rect 132723 79928 132789 79933
rect 132956 79932 133004 79962
rect 130254 79872 132602 79901
rect 130193 79870 132602 79872
rect 132723 79872 132728 79928
rect 132784 79872 132789 79928
rect 130193 79867 130259 79870
rect 132723 79867 132789 79872
rect 132902 79868 132908 79932
rect 132972 79906 133004 79932
rect 133060 79906 133065 79962
rect 134842 79933 134902 80006
rect 139350 79967 139410 80142
rect 145414 80004 145420 80068
rect 145484 80066 145490 80068
rect 145484 80006 146218 80066
rect 145484 80004 145490 80006
rect 135023 79964 135089 79967
rect 134980 79962 135089 79964
rect 132972 79901 133065 79906
rect 133919 79930 133985 79933
rect 134558 79930 134564 79932
rect 133919 79928 134564 79930
rect 132972 79870 133016 79901
rect 133919 79872 133924 79928
rect 133980 79872 134564 79928
rect 133919 79870 134564 79872
rect 132972 79868 132978 79870
rect 133919 79867 133985 79870
rect 134558 79868 134564 79870
rect 134628 79868 134634 79932
rect 134839 79928 134905 79933
rect 134839 79872 134844 79928
rect 134900 79872 134905 79928
rect 134839 79867 134905 79872
rect 134980 79906 135028 79962
rect 135084 79906 135089 79962
rect 134980 79901 135089 79906
rect 135391 79964 135457 79967
rect 135391 79962 135500 79964
rect 135391 79906 135396 79962
rect 135452 79930 135500 79962
rect 136403 79962 136469 79967
rect 135846 79930 135852 79932
rect 135452 79906 135852 79930
rect 135391 79901 135852 79906
rect 132726 79797 132786 79867
rect 131614 79732 131620 79796
rect 131684 79794 131690 79796
rect 132217 79794 132283 79797
rect 131684 79792 132283 79794
rect 131684 79736 132222 79792
rect 132278 79736 132283 79792
rect 131684 79734 132283 79736
rect 131684 79732 131690 79734
rect 132217 79731 132283 79734
rect 132677 79794 132786 79797
rect 133086 79794 133092 79796
rect 132677 79792 133092 79794
rect 132677 79736 132682 79792
rect 132738 79736 133092 79792
rect 132677 79734 133092 79736
rect 132677 79731 132743 79734
rect 133086 79732 133092 79734
rect 133156 79732 133162 79796
rect 133321 79794 133387 79797
rect 133638 79794 133644 79796
rect 133321 79792 133644 79794
rect 133321 79736 133326 79792
rect 133382 79736 133644 79792
rect 133321 79734 133644 79736
rect 133321 79731 133387 79734
rect 133638 79732 133644 79734
rect 133708 79732 133714 79796
rect 134517 79792 134583 79797
rect 134517 79736 134522 79792
rect 134578 79736 134583 79792
rect 134517 79731 134583 79736
rect 134742 79732 134748 79796
rect 134812 79794 134818 79796
rect 134980 79794 135040 79901
rect 135440 79870 135852 79901
rect 135846 79868 135852 79870
rect 135916 79868 135922 79932
rect 136403 79906 136408 79962
rect 136464 79906 136469 79962
rect 136403 79901 136469 79906
rect 136771 79962 136837 79967
rect 136771 79906 136776 79962
rect 136832 79906 136837 79962
rect 136771 79901 136837 79906
rect 137047 79964 137113 79967
rect 137047 79962 137156 79964
rect 137047 79906 137052 79962
rect 137108 79932 137156 79962
rect 138335 79962 138401 79967
rect 137108 79906 137140 79932
rect 137047 79901 137140 79906
rect 135115 79826 135181 79831
rect 135115 79796 135120 79826
rect 135176 79796 135181 79826
rect 134812 79734 135040 79794
rect 134812 79732 134818 79734
rect 135110 79732 135116 79796
rect 135180 79794 135186 79796
rect 135253 79794 135319 79797
rect 135180 79792 135319 79794
rect 135180 79736 135258 79792
rect 135314 79736 135319 79792
rect 135180 79734 135319 79736
rect 135180 79732 135186 79734
rect 135253 79731 135319 79734
rect 132125 79658 132191 79661
rect 133270 79658 133276 79660
rect 132125 79656 133276 79658
rect 132125 79600 132130 79656
rect 132186 79600 133276 79656
rect 132125 79598 133276 79600
rect 132125 79595 132191 79598
rect 133270 79596 133276 79598
rect 133340 79596 133346 79660
rect 134190 79596 134196 79660
rect 134260 79658 134266 79660
rect 134520 79658 134580 79731
rect 136406 79661 136466 79901
rect 136774 79794 136834 79901
rect 137096 79870 137140 79901
rect 137134 79868 137140 79870
rect 137204 79868 137210 79932
rect 137323 79930 137389 79933
rect 137502 79930 137508 79932
rect 137323 79928 137508 79930
rect 137323 79872 137328 79928
rect 137384 79872 137508 79928
rect 137323 79870 137508 79872
rect 137323 79867 137389 79870
rect 137502 79868 137508 79870
rect 137572 79868 137578 79932
rect 137686 79868 137692 79932
rect 137756 79930 137762 79932
rect 137875 79930 137941 79933
rect 138335 79930 138340 79962
rect 137756 79928 137941 79930
rect 137756 79872 137880 79928
rect 137936 79872 137941 79928
rect 137756 79870 137941 79872
rect 137756 79868 137762 79870
rect 137875 79867 137941 79870
rect 138108 79906 138340 79930
rect 138396 79906 138401 79962
rect 139347 79962 139413 79967
rect 138108 79901 138401 79906
rect 138703 79930 138769 79933
rect 138974 79930 138980 79932
rect 138703 79928 138980 79930
rect 138108 79870 138398 79901
rect 138703 79872 138708 79928
rect 138764 79872 138980 79928
rect 138703 79870 138980 79872
rect 136950 79794 136956 79796
rect 136774 79734 136956 79794
rect 136950 79732 136956 79734
rect 137020 79732 137026 79796
rect 137093 79794 137159 79797
rect 137318 79794 137324 79796
rect 137093 79792 137324 79794
rect 137093 79736 137098 79792
rect 137154 79736 137324 79792
rect 137093 79734 137324 79736
rect 137093 79731 137159 79734
rect 137318 79732 137324 79734
rect 137388 79732 137394 79796
rect 134260 79598 134580 79658
rect 134260 79596 134266 79598
rect 134926 79596 134932 79660
rect 134996 79658 135002 79660
rect 135069 79658 135135 79661
rect 134996 79656 135135 79658
rect 134996 79600 135074 79656
rect 135130 79600 135135 79656
rect 134996 79598 135135 79600
rect 134996 79596 135002 79598
rect 135069 79595 135135 79598
rect 135713 79658 135779 79661
rect 136214 79658 136220 79660
rect 135713 79656 136220 79658
rect 135713 79600 135718 79656
rect 135774 79600 136220 79656
rect 135713 79598 136220 79600
rect 135713 79595 135779 79598
rect 136214 79596 136220 79598
rect 136284 79596 136290 79660
rect 136357 79656 136466 79661
rect 136357 79600 136362 79656
rect 136418 79600 136466 79656
rect 136357 79598 136466 79600
rect 136357 79595 136423 79598
rect 136582 79596 136588 79660
rect 136652 79658 136658 79660
rect 137645 79658 137711 79661
rect 136652 79656 137711 79658
rect 136652 79600 137650 79656
rect 137706 79600 137711 79656
rect 136652 79598 137711 79600
rect 138108 79658 138168 79870
rect 138703 79867 138769 79870
rect 138974 79868 138980 79870
rect 139044 79868 139050 79932
rect 139347 79906 139352 79962
rect 139408 79906 139413 79962
rect 142475 79962 142541 79967
rect 144775 79964 144841 79967
rect 139531 79932 139597 79933
rect 139347 79901 139413 79906
rect 139526 79868 139532 79932
rect 139596 79930 139602 79932
rect 139596 79870 139688 79930
rect 139807 79928 139873 79933
rect 139807 79872 139812 79928
rect 139868 79872 139873 79928
rect 140635 79928 140701 79933
rect 139596 79868 139602 79870
rect 139531 79867 139597 79868
rect 139807 79867 139873 79872
rect 140083 79894 140149 79899
rect 138289 79794 138355 79797
rect 138790 79794 138796 79796
rect 138289 79792 138796 79794
rect 138289 79736 138294 79792
rect 138350 79736 138796 79792
rect 138289 79734 138796 79736
rect 138289 79731 138355 79734
rect 138790 79732 138796 79734
rect 138860 79732 138866 79796
rect 139342 79732 139348 79796
rect 139412 79794 139418 79796
rect 139810 79794 139870 79867
rect 140083 79838 140088 79894
rect 140144 79838 140149 79894
rect 140635 79872 140640 79928
rect 140696 79872 140701 79928
rect 140635 79867 140701 79872
rect 140819 79928 140885 79933
rect 140819 79872 140824 79928
rect 140880 79872 140885 79928
rect 140819 79867 140885 79872
rect 140998 79868 141004 79932
rect 141068 79930 141074 79932
rect 141739 79930 141805 79933
rect 141068 79928 141805 79930
rect 141068 79872 141744 79928
rect 141800 79872 141805 79928
rect 142475 79906 142480 79962
rect 142536 79906 142541 79962
rect 144732 79962 144841 79964
rect 142475 79901 142541 79906
rect 141068 79870 141805 79872
rect 141068 79868 141074 79870
rect 141739 79867 141805 79870
rect 140083 79833 140149 79838
rect 139412 79734 139870 79794
rect 139412 79732 139418 79734
rect 138422 79658 138428 79660
rect 138108 79598 138428 79658
rect 136652 79596 136658 79598
rect 137645 79595 137711 79598
rect 138422 79596 138428 79598
rect 138492 79596 138498 79660
rect 138606 79596 138612 79660
rect 138676 79658 138682 79660
rect 139025 79658 139091 79661
rect 139209 79660 139275 79661
rect 138676 79656 139091 79658
rect 138676 79600 139030 79656
rect 139086 79600 139091 79656
rect 138676 79598 139091 79600
rect 138676 79596 138682 79598
rect 139025 79595 139091 79598
rect 139158 79596 139164 79660
rect 139228 79658 139275 79660
rect 139669 79660 139735 79661
rect 139228 79656 139320 79658
rect 139270 79600 139320 79656
rect 139228 79598 139320 79600
rect 139669 79656 139716 79660
rect 139780 79658 139786 79660
rect 140086 79658 140146 79833
rect 140262 79732 140268 79796
rect 140332 79794 140338 79796
rect 140638 79794 140698 79867
rect 140332 79734 140698 79794
rect 140822 79794 140882 79867
rect 142478 79797 142538 79901
rect 142843 79894 142909 79899
rect 142843 79838 142848 79894
rect 142904 79838 142909 79894
rect 143022 79868 143028 79932
rect 143092 79930 143098 79932
rect 143303 79930 143369 79933
rect 143092 79928 143369 79930
rect 143092 79872 143308 79928
rect 143364 79872 143369 79928
rect 143092 79870 143369 79872
rect 143092 79868 143098 79870
rect 143303 79867 143369 79870
rect 143487 79928 143553 79933
rect 143487 79872 143492 79928
rect 143548 79872 143553 79928
rect 143487 79867 143553 79872
rect 143763 79928 143829 79933
rect 143763 79872 143768 79928
rect 143824 79872 143829 79928
rect 143763 79867 143829 79872
rect 144310 79868 144316 79932
rect 144380 79930 144386 79932
rect 144732 79930 144780 79962
rect 144380 79906 144780 79930
rect 144836 79906 144841 79962
rect 145235 79962 145301 79967
rect 144380 79901 144841 79906
rect 144380 79870 144792 79901
rect 144380 79868 144386 79870
rect 145046 79868 145052 79932
rect 145116 79930 145122 79932
rect 145235 79930 145240 79962
rect 145116 79906 145240 79930
rect 145296 79906 145301 79962
rect 146158 79933 146218 80006
rect 145116 79901 145301 79906
rect 145116 79870 145298 79901
rect 145116 79868 145122 79870
rect 145414 79868 145420 79932
rect 145484 79930 145490 79932
rect 145603 79930 145669 79933
rect 145484 79928 145669 79930
rect 145484 79872 145608 79928
rect 145664 79872 145669 79928
rect 145484 79870 145669 79872
rect 145484 79868 145490 79870
rect 145603 79867 145669 79870
rect 145971 79928 146037 79933
rect 146155 79930 146221 79933
rect 145971 79872 145976 79928
rect 146032 79872 146037 79928
rect 145971 79867 146037 79872
rect 146112 79928 146221 79930
rect 146112 79872 146160 79928
rect 146216 79872 146221 79928
rect 146112 79867 146221 79872
rect 146296 79930 146356 80278
rect 147814 80202 147874 80550
rect 164182 80548 164188 80612
rect 164252 80610 164258 80612
rect 172470 80610 172530 80686
rect 176326 80610 176332 80612
rect 164252 80550 168850 80610
rect 172470 80550 176332 80610
rect 164252 80548 164258 80550
rect 161238 80412 161244 80476
rect 161308 80474 161314 80476
rect 168790 80474 168850 80550
rect 176326 80548 176332 80550
rect 176396 80548 176402 80612
rect 177576 80610 177636 80822
rect 179324 80880 523191 80882
rect 179324 80824 199106 80880
rect 199162 80824 523130 80880
rect 523186 80824 523191 80880
rect 179324 80822 523191 80824
rect 179324 80749 179384 80822
rect 199101 80819 199167 80822
rect 523125 80819 523191 80822
rect 179321 80744 179387 80749
rect 179321 80688 179326 80744
rect 179382 80688 179387 80744
rect 179321 80683 179387 80688
rect 179597 80748 179663 80749
rect 179597 80744 179644 80748
rect 179708 80746 179714 80748
rect 179873 80746 179939 80749
rect 198958 80746 198964 80748
rect 179597 80688 179602 80744
rect 179597 80684 179644 80688
rect 179708 80686 179754 80746
rect 179873 80744 198964 80746
rect 179873 80688 179878 80744
rect 179934 80688 198964 80744
rect 179873 80686 198964 80688
rect 179708 80684 179714 80686
rect 179597 80683 179663 80684
rect 179873 80683 179939 80686
rect 198958 80684 198964 80686
rect 199028 80746 199034 80748
rect 525793 80746 525859 80749
rect 199028 80744 525859 80746
rect 199028 80688 525798 80744
rect 525854 80688 525859 80744
rect 199028 80686 525859 80688
rect 199028 80684 199034 80686
rect 525793 80683 525859 80686
rect 177757 80610 177823 80613
rect 177576 80608 177823 80610
rect 177576 80552 177762 80608
rect 177818 80552 177823 80608
rect 177576 80550 177823 80552
rect 177757 80547 177823 80550
rect 178125 80474 178191 80477
rect 161308 80414 167056 80474
rect 168790 80472 178191 80474
rect 168790 80416 178130 80472
rect 178186 80416 178191 80472
rect 168790 80414 178191 80416
rect 161308 80412 161314 80414
rect 156638 80276 156644 80340
rect 156708 80338 156714 80340
rect 157190 80338 157196 80340
rect 156708 80278 157196 80338
rect 156708 80276 156714 80278
rect 157190 80276 157196 80278
rect 157260 80276 157266 80340
rect 160870 80276 160876 80340
rect 160940 80338 160946 80340
rect 166996 80338 167056 80414
rect 178125 80411 178191 80414
rect 181437 80474 181503 80477
rect 188429 80474 188495 80477
rect 181437 80472 188495 80474
rect 181437 80416 181442 80472
rect 181498 80416 188434 80472
rect 188490 80416 188495 80472
rect 181437 80414 188495 80416
rect 181437 80411 181503 80414
rect 188429 80411 188495 80414
rect 160940 80278 161260 80338
rect 166996 80278 168436 80338
rect 160940 80276 160946 80278
rect 147814 80142 149208 80202
rect 149148 80066 149208 80142
rect 150750 80140 150756 80204
rect 150820 80202 150826 80204
rect 150820 80142 151462 80202
rect 150820 80140 150826 80142
rect 151402 80066 151462 80142
rect 154798 80140 154804 80204
rect 154868 80202 154874 80204
rect 154868 80142 155924 80202
rect 154868 80140 154874 80142
rect 155718 80066 155724 80068
rect 149148 80006 149530 80066
rect 151402 80006 151692 80066
rect 146891 79962 146957 79967
rect 148455 79964 148521 79967
rect 146615 79930 146681 79933
rect 146296 79928 146681 79930
rect 146296 79872 146620 79928
rect 146676 79872 146681 79928
rect 146891 79906 146896 79962
rect 146952 79906 146957 79962
rect 148412 79962 148521 79964
rect 146891 79901 146957 79906
rect 147259 79930 147325 79933
rect 148412 79930 148460 79962
rect 147259 79928 147460 79930
rect 146296 79870 146681 79872
rect 142843 79833 142909 79838
rect 140998 79794 141004 79796
rect 140822 79734 141004 79794
rect 140332 79732 140338 79734
rect 140998 79732 141004 79734
rect 141068 79732 141074 79796
rect 141187 79794 141253 79797
rect 141550 79794 141556 79796
rect 141187 79792 141556 79794
rect 141187 79736 141192 79792
rect 141248 79736 141556 79792
rect 141187 79734 141556 79736
rect 141187 79731 141253 79734
rect 141550 79732 141556 79734
rect 141620 79732 141626 79796
rect 141923 79792 141989 79797
rect 142199 79794 142265 79797
rect 141923 79736 141928 79792
rect 141984 79736 141989 79792
rect 141923 79731 141989 79736
rect 142064 79792 142265 79794
rect 142064 79736 142204 79792
rect 142260 79736 142265 79792
rect 142064 79734 142265 79736
rect 142478 79792 142587 79797
rect 142478 79736 142526 79792
rect 142582 79736 142587 79792
rect 142478 79734 142587 79736
rect 140630 79658 140636 79660
rect 139669 79600 139674 79656
rect 139228 79596 139275 79598
rect 139209 79595 139275 79596
rect 139669 79596 139716 79600
rect 139780 79598 139826 79658
rect 140086 79598 140636 79658
rect 139780 79596 139786 79598
rect 140630 79596 140636 79598
rect 140700 79596 140706 79660
rect 140773 79658 140839 79661
rect 141190 79658 141250 79731
rect 141417 79660 141483 79661
rect 140773 79656 141250 79658
rect 140773 79600 140778 79656
rect 140834 79600 141250 79656
rect 140773 79598 141250 79600
rect 139669 79595 139735 79596
rect 140773 79595 140839 79598
rect 141366 79596 141372 79660
rect 141436 79658 141483 79660
rect 141693 79658 141759 79661
rect 141926 79658 141986 79731
rect 141436 79656 141528 79658
rect 141478 79600 141528 79656
rect 141436 79598 141528 79600
rect 141693 79656 141986 79658
rect 141693 79600 141698 79656
rect 141754 79600 141986 79656
rect 141693 79598 141986 79600
rect 142064 79658 142124 79734
rect 142199 79731 142265 79734
rect 142521 79731 142587 79734
rect 142429 79658 142495 79661
rect 142064 79656 142495 79658
rect 142064 79600 142434 79656
rect 142490 79600 142495 79656
rect 142064 79598 142495 79600
rect 141436 79596 141483 79598
rect 141417 79595 141483 79596
rect 141693 79595 141759 79598
rect 142429 79595 142495 79598
rect 142613 79658 142679 79661
rect 142846 79658 142906 79833
rect 142613 79656 142906 79658
rect 142613 79600 142618 79656
rect 142674 79600 142906 79656
rect 142613 79598 142906 79600
rect 143490 79661 143550 79867
rect 143490 79656 143599 79661
rect 143490 79600 143538 79656
rect 143594 79600 143599 79656
rect 143490 79598 143599 79600
rect 143766 79658 143826 79867
rect 145974 79797 146034 79867
rect 146112 79797 146172 79867
rect 144494 79732 144500 79796
rect 144564 79794 144570 79796
rect 144683 79794 144749 79797
rect 144564 79792 144749 79794
rect 144564 79736 144688 79792
rect 144744 79736 144749 79792
rect 144564 79734 144749 79736
rect 144564 79732 144570 79734
rect 144683 79731 144749 79734
rect 144862 79732 144868 79796
rect 144932 79794 144938 79796
rect 145741 79794 145807 79797
rect 144932 79792 145807 79794
rect 144932 79736 145746 79792
rect 145802 79736 145807 79792
rect 144932 79734 145807 79736
rect 144932 79732 144938 79734
rect 145741 79731 145807 79734
rect 145925 79792 146034 79797
rect 145925 79736 145930 79792
rect 145986 79736 146034 79792
rect 145925 79734 146034 79736
rect 146109 79792 146175 79797
rect 146109 79736 146114 79792
rect 146170 79736 146175 79792
rect 145925 79731 145991 79734
rect 146109 79731 146175 79736
rect 144361 79658 144427 79661
rect 143766 79656 144427 79658
rect 143766 79600 144366 79656
rect 144422 79600 144427 79656
rect 143766 79598 144427 79600
rect 146296 79658 146356 79870
rect 146615 79867 146681 79870
rect 146894 79797 146954 79901
rect 147259 79872 147264 79928
rect 147320 79872 147460 79928
rect 147259 79870 147460 79872
rect 147259 79867 147325 79870
rect 146894 79792 147003 79797
rect 146894 79736 146942 79792
rect 146998 79736 147003 79792
rect 146894 79734 147003 79736
rect 146937 79731 147003 79734
rect 146477 79658 146543 79661
rect 146296 79656 146543 79658
rect 146296 79600 146482 79656
rect 146538 79600 146543 79656
rect 146296 79598 146543 79600
rect 142613 79595 142679 79598
rect 143533 79595 143599 79598
rect 144361 79595 144427 79598
rect 146477 79595 146543 79598
rect 146886 79596 146892 79660
rect 146956 79658 146962 79660
rect 147400 79658 147460 79870
rect 148228 79906 148460 79930
rect 148516 79906 148521 79962
rect 148639 79964 148705 79967
rect 148639 79962 148716 79964
rect 148639 79932 148644 79962
rect 148228 79901 148521 79906
rect 148228 79870 148472 79901
rect 148228 79797 148288 79870
rect 148588 79868 148594 79932
rect 148700 79906 148716 79962
rect 148658 79904 148716 79906
rect 148915 79928 148981 79933
rect 148658 79901 148705 79904
rect 148658 79870 148702 79901
rect 148915 79872 148920 79928
rect 148976 79872 148981 79928
rect 148658 79868 148664 79870
rect 148915 79867 148981 79872
rect 149099 79930 149165 79933
rect 149099 79928 149346 79930
rect 149099 79872 149104 79928
rect 149160 79872 149346 79928
rect 149099 79870 149346 79872
rect 149099 79867 149165 79870
rect 148041 79796 148107 79797
rect 147990 79732 147996 79796
rect 148060 79794 148107 79796
rect 148060 79792 148152 79794
rect 148102 79736 148152 79792
rect 148060 79734 148152 79736
rect 148225 79792 148291 79797
rect 148225 79736 148230 79792
rect 148286 79736 148291 79792
rect 148060 79732 148107 79734
rect 148041 79731 148107 79732
rect 148225 79731 148291 79736
rect 148358 79732 148364 79796
rect 148428 79794 148434 79796
rect 148918 79794 148978 79867
rect 149094 79794 149100 79796
rect 148428 79734 149100 79794
rect 148428 79732 148434 79734
rect 149094 79732 149100 79734
rect 149164 79732 149170 79796
rect 149286 79661 149346 79870
rect 147581 79658 147647 79661
rect 146956 79656 147647 79658
rect 146956 79600 147586 79656
rect 147642 79600 147647 79656
rect 146956 79598 147647 79600
rect 146956 79596 146962 79598
rect 147581 79595 147647 79598
rect 149237 79656 149346 79661
rect 149237 79600 149242 79656
rect 149298 79600 149346 79656
rect 149237 79598 149346 79600
rect 149470 79658 149530 80006
rect 151632 79967 151692 80006
rect 154990 80006 155724 80066
rect 150847 79964 150913 79967
rect 150847 79962 150956 79964
rect 150203 79932 150269 79933
rect 150387 79932 150453 79933
rect 150198 79930 150204 79932
rect 150112 79870 150204 79930
rect 150198 79868 150204 79870
rect 150268 79868 150274 79932
rect 150382 79868 150388 79932
rect 150452 79930 150458 79932
rect 150452 79870 150544 79930
rect 150847 79906 150852 79962
rect 150908 79932 150956 79962
rect 151632 79962 151741 79967
rect 150908 79906 150940 79932
rect 150847 79901 150940 79906
rect 150452 79868 150458 79870
rect 150896 79868 150940 79901
rect 151004 79868 151010 79932
rect 151123 79930 151189 79933
rect 151486 79930 151492 79932
rect 151123 79928 151492 79930
rect 151123 79872 151128 79928
rect 151184 79872 151492 79928
rect 151123 79870 151492 79872
rect 150203 79867 150269 79868
rect 150387 79867 150453 79868
rect 150896 79797 150956 79868
rect 151123 79867 151189 79870
rect 151486 79868 151492 79870
rect 151556 79868 151562 79932
rect 151632 79906 151680 79962
rect 151736 79906 151741 79962
rect 151632 79904 151741 79906
rect 151675 79901 151741 79904
rect 151859 79962 151925 79967
rect 151859 79906 151864 79962
rect 151920 79906 151925 79962
rect 154990 79933 155050 80006
rect 155718 80004 155724 80006
rect 155788 80004 155794 80068
rect 155864 79933 155924 80142
rect 159582 80140 159588 80204
rect 159652 80202 159658 80204
rect 159652 80142 159972 80202
rect 159652 80140 159658 80142
rect 156270 80004 156276 80068
rect 156340 80066 156346 80068
rect 156340 80006 158776 80066
rect 156340 80004 156346 80006
rect 153883 79932 153949 79933
rect 151859 79901 151925 79906
rect 149646 79732 149652 79796
rect 149716 79794 149722 79796
rect 150249 79794 150315 79797
rect 149716 79792 150315 79794
rect 149716 79736 150254 79792
rect 150310 79736 150315 79792
rect 149716 79734 150315 79736
rect 149716 79732 149722 79734
rect 150249 79731 150315 79734
rect 150893 79792 150959 79797
rect 150893 79736 150898 79792
rect 150954 79736 150959 79792
rect 150893 79731 150959 79736
rect 151031 79794 151097 79797
rect 151031 79792 151140 79794
rect 151031 79736 151036 79792
rect 151092 79736 151140 79792
rect 151031 79731 151140 79736
rect 151080 79661 151140 79731
rect 151862 79661 151922 79901
rect 152222 79868 152228 79932
rect 152292 79930 152298 79932
rect 152292 79899 152566 79930
rect 152292 79894 152569 79899
rect 152292 79870 152508 79894
rect 152292 79868 152298 79870
rect 152503 79838 152508 79870
rect 152564 79838 152569 79894
rect 153878 79868 153884 79932
rect 153948 79930 153954 79932
rect 153948 79870 154040 79930
rect 154435 79928 154501 79933
rect 154435 79872 154440 79928
rect 154496 79872 154501 79928
rect 153948 79868 153954 79870
rect 153883 79867 153949 79868
rect 154435 79867 154501 79872
rect 154987 79928 155053 79933
rect 154987 79872 154992 79928
rect 155048 79872 155053 79928
rect 154987 79867 155053 79872
rect 155350 79868 155356 79932
rect 155420 79930 155426 79932
rect 155539 79930 155605 79933
rect 155420 79928 155648 79930
rect 155420 79872 155544 79928
rect 155600 79872 155648 79928
rect 155420 79870 155648 79872
rect 155420 79868 155426 79870
rect 155539 79867 155648 79870
rect 155815 79928 155924 79933
rect 155815 79872 155820 79928
rect 155876 79872 155924 79928
rect 155815 79870 155924 79872
rect 155815 79867 155881 79870
rect 156454 79868 156460 79932
rect 156524 79930 156530 79932
rect 157011 79930 157077 79933
rect 157195 79932 157261 79933
rect 156524 79928 157077 79930
rect 156524 79872 157016 79928
rect 157072 79872 157077 79928
rect 156524 79870 157077 79872
rect 156524 79868 156530 79870
rect 157011 79867 157077 79870
rect 157190 79868 157196 79932
rect 157260 79930 157266 79932
rect 157747 79930 157813 79933
rect 157926 79930 157932 79932
rect 157260 79870 157352 79930
rect 157704 79928 157932 79930
rect 157704 79872 157752 79928
rect 157808 79872 157932 79928
rect 157704 79870 157932 79872
rect 157260 79868 157266 79870
rect 157195 79867 157261 79868
rect 157704 79867 157813 79870
rect 157926 79868 157932 79870
rect 157996 79868 158002 79932
rect 158294 79868 158300 79932
rect 158364 79930 158370 79932
rect 158575 79930 158641 79933
rect 158364 79928 158641 79930
rect 158364 79872 158580 79928
rect 158636 79872 158641 79928
rect 158364 79870 158641 79872
rect 158364 79868 158370 79870
rect 158575 79867 158641 79870
rect 152503 79833 152569 79838
rect 152227 79796 152293 79797
rect 152222 79794 152228 79796
rect 152136 79734 152228 79794
rect 152222 79732 152228 79734
rect 152292 79732 152298 79796
rect 152227 79731 152293 79732
rect 149697 79658 149763 79661
rect 149470 79656 149763 79658
rect 149470 79600 149702 79656
rect 149758 79600 149763 79656
rect 149470 79598 149763 79600
rect 149237 79595 149303 79598
rect 149697 79595 149763 79598
rect 149830 79596 149836 79660
rect 149900 79658 149906 79660
rect 150525 79658 150591 79661
rect 151077 79658 151143 79661
rect 149900 79656 150591 79658
rect 149900 79600 150530 79656
rect 150586 79600 150591 79656
rect 149900 79598 150591 79600
rect 149900 79596 149906 79598
rect 150525 79595 150591 79598
rect 150942 79656 151143 79658
rect 150942 79600 151082 79656
rect 151138 79600 151143 79656
rect 150942 79598 151143 79600
rect 117957 79522 118023 79525
rect 150942 79522 151002 79598
rect 151077 79595 151143 79598
rect 151261 79660 151327 79661
rect 151261 79656 151308 79660
rect 151372 79658 151378 79660
rect 151261 79600 151266 79656
rect 151261 79596 151308 79600
rect 151372 79598 151418 79658
rect 151862 79656 151971 79661
rect 151862 79600 151910 79656
rect 151966 79600 151971 79656
rect 151862 79598 151971 79600
rect 152506 79658 152566 79833
rect 153510 79794 153516 79796
rect 153472 79732 153516 79794
rect 153580 79794 153586 79796
rect 154438 79794 154498 79867
rect 153580 79734 154498 79794
rect 154573 79794 154639 79797
rect 155217 79794 155283 79797
rect 155350 79794 155356 79796
rect 154573 79792 155356 79794
rect 154573 79736 154578 79792
rect 154634 79736 155222 79792
rect 155278 79736 155356 79792
rect 154573 79734 155356 79736
rect 153580 79732 153586 79734
rect 152641 79658 152707 79661
rect 152506 79656 152707 79658
rect 152506 79600 152646 79656
rect 152702 79600 152707 79656
rect 152506 79598 152707 79600
rect 151372 79596 151378 79598
rect 151261 79595 151327 79596
rect 151905 79595 151971 79598
rect 152641 79595 152707 79598
rect 153472 79525 153532 79732
rect 154573 79731 154639 79734
rect 155217 79731 155283 79734
rect 155350 79732 155356 79734
rect 155420 79732 155426 79796
rect 155588 79661 155648 79867
rect 157704 79797 157764 79867
rect 156367 79792 156433 79797
rect 156367 79736 156372 79792
rect 156428 79736 156433 79792
rect 156367 79731 156433 79736
rect 156643 79794 156709 79797
rect 157006 79794 157012 79796
rect 156643 79792 157012 79794
rect 156643 79736 156648 79792
rect 156704 79736 157012 79792
rect 156643 79734 157012 79736
rect 156643 79731 156709 79734
rect 157006 79732 157012 79734
rect 157076 79732 157082 79796
rect 157701 79792 157767 79797
rect 157701 79736 157706 79792
rect 157762 79736 157767 79792
rect 157701 79731 157767 79736
rect 158716 79794 158776 80006
rect 159912 79967 159972 80142
rect 159495 79962 159561 79967
rect 158846 79868 158852 79932
rect 158916 79930 158922 79932
rect 159495 79930 159500 79962
rect 158916 79906 159500 79930
rect 159556 79906 159561 79962
rect 159912 79962 160021 79967
rect 159679 79930 159745 79933
rect 158916 79901 159561 79906
rect 159636 79928 159745 79930
rect 158916 79870 159558 79901
rect 159636 79872 159684 79928
rect 159740 79872 159745 79928
rect 159912 79906 159960 79962
rect 160016 79906 160021 79962
rect 160323 79932 160389 79933
rect 160318 79930 160324 79932
rect 159912 79904 160021 79906
rect 159955 79901 160021 79904
rect 158916 79868 158922 79870
rect 159636 79867 159745 79872
rect 160232 79870 160324 79930
rect 160318 79868 160324 79870
rect 160388 79868 160394 79932
rect 160323 79867 160389 79868
rect 158851 79794 158917 79797
rect 158716 79792 158917 79794
rect 158716 79736 158856 79792
rect 158912 79736 158917 79792
rect 158716 79734 158917 79736
rect 158851 79731 158917 79734
rect 159030 79732 159036 79796
rect 159100 79794 159106 79796
rect 159403 79794 159469 79797
rect 159100 79792 159469 79794
rect 159100 79736 159408 79792
rect 159464 79736 159469 79792
rect 159100 79734 159469 79736
rect 159100 79732 159106 79734
rect 159403 79731 159469 79734
rect 153745 79658 153811 79661
rect 154205 79660 154271 79661
rect 154062 79658 154068 79660
rect 153745 79656 154068 79658
rect 153745 79600 153750 79656
rect 153806 79600 154068 79656
rect 153745 79598 154068 79600
rect 153745 79595 153811 79598
rect 154062 79596 154068 79598
rect 154132 79596 154138 79660
rect 154205 79656 154252 79660
rect 154316 79658 154322 79660
rect 154205 79600 154210 79656
rect 154205 79596 154252 79600
rect 154316 79598 154362 79658
rect 155585 79656 155651 79661
rect 155585 79600 155590 79656
rect 155646 79600 155651 79656
rect 154316 79596 154322 79598
rect 154205 79595 154271 79596
rect 155585 79595 155651 79600
rect 117957 79520 151002 79522
rect 117957 79464 117962 79520
rect 118018 79464 151002 79520
rect 117957 79462 151002 79464
rect 117957 79459 118023 79462
rect 152590 79460 152596 79524
rect 152660 79522 152666 79524
rect 152733 79522 152799 79525
rect 152660 79520 152799 79522
rect 152660 79464 152738 79520
rect 152794 79464 152799 79520
rect 152660 79462 152799 79464
rect 152660 79460 152666 79462
rect 152733 79459 152799 79462
rect 153469 79520 153535 79525
rect 153469 79464 153474 79520
rect 153530 79464 153535 79520
rect 153469 79459 153535 79464
rect 153694 79460 153700 79524
rect 153764 79522 153770 79524
rect 154297 79522 154363 79525
rect 155769 79524 155835 79525
rect 153764 79520 154363 79522
rect 153764 79464 154302 79520
rect 154358 79464 154363 79520
rect 153764 79462 154363 79464
rect 153764 79460 153770 79462
rect 154297 79459 154363 79462
rect 155718 79460 155724 79524
rect 155788 79522 155835 79524
rect 155788 79520 155880 79522
rect 155830 79464 155880 79520
rect 155788 79462 155880 79464
rect 155788 79460 155835 79462
rect 155769 79459 155835 79460
rect 124121 79386 124187 79389
rect 130101 79386 130167 79389
rect 124121 79384 130167 79386
rect 124121 79328 124126 79384
rect 124182 79328 130106 79384
rect 130162 79328 130167 79384
rect 124121 79326 130167 79328
rect 124121 79323 124187 79326
rect 130101 79323 130167 79326
rect 131982 79324 131988 79388
rect 132052 79386 132058 79388
rect 150801 79386 150867 79389
rect 151445 79386 151511 79389
rect 132052 79384 151511 79386
rect 132052 79328 150806 79384
rect 150862 79328 151450 79384
rect 151506 79328 151511 79384
rect 132052 79326 151511 79328
rect 132052 79324 132058 79326
rect 150801 79323 150867 79326
rect 151445 79323 151511 79326
rect 152181 79386 152247 79389
rect 152774 79386 152780 79388
rect 152181 79384 152780 79386
rect 152181 79328 152186 79384
rect 152242 79328 152780 79384
rect 152181 79326 152780 79328
rect 152181 79323 152247 79326
rect 152774 79324 152780 79326
rect 152844 79324 152850 79388
rect 153878 79324 153884 79388
rect 153948 79386 153954 79388
rect 154205 79386 154271 79389
rect 153948 79384 154271 79386
rect 153948 79328 154210 79384
rect 154266 79328 154271 79384
rect 153948 79326 154271 79328
rect 156370 79386 156430 79731
rect 159636 79661 159696 79867
rect 161200 79797 161260 80278
rect 167310 80140 167316 80204
rect 167380 80202 167386 80204
rect 168376 80202 168436 80278
rect 170622 80276 170628 80340
rect 170692 80338 170698 80340
rect 170692 80278 186330 80338
rect 170692 80276 170698 80278
rect 170254 80202 170260 80204
rect 167380 80142 168298 80202
rect 168376 80142 168482 80202
rect 167380 80140 167386 80142
rect 161974 80004 161980 80068
rect 162044 80066 162050 80068
rect 165470 80066 165476 80068
rect 162044 80006 162778 80066
rect 162044 80004 162050 80006
rect 162718 79933 162778 80006
rect 165110 80006 165476 80066
rect 162899 79962 162965 79967
rect 161427 79932 161493 79933
rect 161422 79868 161428 79932
rect 161492 79930 161498 79932
rect 161703 79930 161769 79933
rect 161492 79870 161584 79930
rect 161703 79928 161904 79930
rect 161703 79872 161708 79928
rect 161764 79872 161904 79928
rect 161703 79870 161904 79872
rect 161492 79868 161498 79870
rect 161427 79867 161493 79868
rect 161703 79867 161769 79870
rect 160231 79794 160297 79797
rect 160737 79796 160803 79797
rect 160188 79792 160297 79794
rect 160188 79736 160236 79792
rect 160292 79736 160297 79792
rect 160188 79731 160297 79736
rect 160686 79732 160692 79796
rect 160756 79794 160803 79796
rect 160756 79792 160848 79794
rect 160798 79736 160848 79792
rect 160756 79734 160848 79736
rect 161197 79792 161263 79797
rect 161197 79736 161202 79792
rect 161258 79736 161263 79792
rect 160756 79732 160803 79734
rect 160737 79731 160803 79732
rect 161197 79731 161263 79736
rect 156822 79596 156828 79660
rect 156892 79658 156898 79660
rect 156965 79658 157031 79661
rect 157793 79660 157859 79661
rect 157742 79658 157748 79660
rect 156892 79656 157031 79658
rect 156892 79600 156970 79656
rect 157026 79600 157031 79656
rect 156892 79598 157031 79600
rect 157702 79598 157748 79658
rect 157812 79656 157859 79660
rect 158069 79660 158135 79661
rect 158069 79658 158116 79660
rect 157854 79600 157859 79656
rect 156892 79596 156898 79598
rect 156965 79595 157031 79598
rect 157742 79596 157748 79598
rect 157812 79596 157859 79600
rect 158024 79656 158116 79658
rect 158024 79600 158074 79656
rect 158024 79598 158116 79600
rect 157793 79595 157859 79596
rect 158069 79596 158116 79598
rect 158180 79596 158186 79660
rect 158662 79596 158668 79660
rect 158732 79658 158738 79660
rect 159633 79658 159699 79661
rect 160188 79658 160248 79731
rect 160921 79660 160987 79661
rect 158732 79656 159699 79658
rect 158732 79600 159638 79656
rect 159694 79600 159699 79656
rect 158732 79598 159699 79600
rect 158732 79596 158738 79598
rect 158069 79595 158135 79596
rect 159633 79595 159699 79598
rect 159774 79598 160248 79658
rect 157558 79460 157564 79524
rect 157628 79522 157634 79524
rect 157793 79522 157859 79525
rect 157628 79520 157859 79522
rect 157628 79464 157798 79520
rect 157854 79464 157859 79520
rect 157628 79462 157859 79464
rect 157628 79460 157634 79462
rect 157793 79459 157859 79462
rect 156822 79386 156828 79388
rect 156370 79326 156828 79386
rect 153948 79324 153954 79326
rect 154205 79323 154271 79326
rect 156822 79324 156828 79326
rect 156892 79324 156898 79388
rect 125358 79188 125364 79252
rect 125428 79250 125434 79252
rect 144821 79250 144887 79253
rect 125428 79248 144887 79250
rect 125428 79192 144826 79248
rect 144882 79192 144887 79248
rect 125428 79190 144887 79192
rect 125428 79188 125434 79190
rect 144821 79187 144887 79190
rect 145230 79188 145236 79252
rect 145300 79250 145306 79252
rect 147121 79250 147187 79253
rect 145300 79248 147187 79250
rect 145300 79192 147126 79248
rect 147182 79192 147187 79248
rect 145300 79190 147187 79192
rect 145300 79188 145306 79190
rect 147121 79187 147187 79190
rect 148726 79188 148732 79252
rect 148796 79250 148802 79252
rect 158713 79250 158779 79253
rect 159081 79250 159147 79253
rect 148796 79248 159147 79250
rect 148796 79192 158718 79248
rect 158774 79192 159086 79248
rect 159142 79192 159147 79248
rect 148796 79190 159147 79192
rect 148796 79188 148802 79190
rect 158713 79187 158779 79190
rect 159081 79187 159147 79190
rect 126646 79052 126652 79116
rect 126716 79114 126722 79116
rect 138054 79114 138060 79116
rect 126716 79054 138060 79114
rect 126716 79052 126722 79054
rect 138054 79052 138060 79054
rect 138124 79052 138130 79116
rect 145414 79114 145420 79116
rect 139350 79054 145420 79114
rect 125174 78916 125180 78980
rect 125244 78978 125250 78980
rect 139350 78978 139410 79054
rect 145414 79052 145420 79054
rect 145484 79052 145490 79116
rect 146702 79052 146708 79116
rect 146772 79114 146778 79116
rect 147070 79114 147076 79116
rect 146772 79054 147076 79114
rect 146772 79052 146778 79054
rect 147070 79052 147076 79054
rect 147140 79114 147146 79116
rect 147489 79114 147555 79117
rect 147140 79112 147555 79114
rect 147140 79056 147494 79112
rect 147550 79056 147555 79112
rect 147140 79054 147555 79056
rect 147140 79052 147146 79054
rect 147489 79051 147555 79054
rect 148174 79052 148180 79116
rect 148244 79114 148250 79116
rect 148961 79114 149027 79117
rect 148244 79112 149027 79114
rect 148244 79056 148966 79112
rect 149022 79056 149027 79112
rect 148244 79054 149027 79056
rect 148244 79052 148250 79054
rect 148961 79051 149027 79054
rect 149145 79114 149211 79117
rect 149830 79114 149836 79116
rect 149145 79112 149836 79114
rect 149145 79056 149150 79112
rect 149206 79056 149836 79112
rect 149145 79054 149836 79056
rect 149145 79051 149211 79054
rect 149830 79052 149836 79054
rect 149900 79052 149906 79116
rect 150014 79052 150020 79116
rect 150084 79114 150090 79116
rect 159774 79114 159834 79598
rect 160870 79596 160876 79660
rect 160940 79658 160987 79660
rect 161844 79658 161904 79870
rect 162158 79868 162164 79932
rect 162228 79930 162234 79932
rect 162439 79930 162505 79933
rect 162228 79928 162505 79930
rect 162228 79872 162444 79928
rect 162500 79872 162505 79928
rect 162228 79870 162505 79872
rect 162228 79868 162234 79870
rect 162439 79867 162505 79870
rect 162715 79928 162781 79933
rect 162715 79872 162720 79928
rect 162776 79872 162781 79928
rect 162899 79906 162904 79962
rect 162960 79906 162965 79962
rect 162899 79901 162965 79906
rect 162715 79867 162781 79872
rect 162442 79661 162502 79867
rect 162718 79661 162778 79867
rect 162902 79797 162962 79901
rect 163446 79868 163452 79932
rect 163516 79930 163522 79932
rect 163911 79930 163977 79933
rect 163516 79928 163977 79930
rect 163516 79872 163916 79928
rect 163972 79872 163977 79928
rect 163516 79870 163977 79872
rect 163516 79868 163522 79870
rect 163911 79867 163977 79870
rect 164371 79928 164437 79933
rect 164371 79872 164376 79928
rect 164432 79872 164437 79928
rect 164371 79867 164437 79872
rect 164739 79930 164805 79933
rect 165110 79930 165170 80006
rect 165470 80004 165476 80006
rect 165540 80004 165546 80068
rect 166390 80066 166396 80068
rect 166030 80006 166396 80066
rect 165659 79962 165725 79967
rect 165291 79932 165357 79933
rect 164739 79928 165170 79930
rect 164739 79872 164744 79928
rect 164800 79872 165170 79928
rect 164739 79870 165170 79872
rect 164739 79867 164805 79870
rect 165286 79868 165292 79932
rect 165356 79930 165362 79932
rect 165356 79870 165448 79930
rect 165659 79906 165664 79962
rect 165720 79906 165725 79962
rect 166030 79933 166090 80006
rect 166390 80004 166396 80006
rect 166460 80004 166466 80068
rect 168238 79967 168298 80142
rect 167775 79964 167841 79967
rect 167732 79962 167841 79964
rect 165659 79901 165725 79906
rect 166027 79928 166093 79933
rect 166579 79932 166645 79933
rect 166947 79932 167013 79933
rect 166574 79930 166580 79932
rect 165356 79868 165362 79870
rect 165291 79867 165357 79868
rect 162853 79792 162962 79797
rect 162853 79736 162858 79792
rect 162914 79736 162962 79792
rect 162853 79734 162962 79736
rect 164374 79797 164434 79867
rect 164374 79792 164483 79797
rect 164374 79736 164422 79792
rect 164478 79736 164483 79792
rect 164374 79734 164483 79736
rect 162853 79731 162919 79734
rect 164417 79731 164483 79734
rect 164693 79796 164759 79797
rect 164693 79792 164740 79796
rect 164804 79794 164810 79796
rect 164923 79794 164989 79797
rect 165102 79794 165108 79796
rect 164693 79736 164698 79792
rect 164693 79732 164740 79736
rect 164804 79734 164850 79794
rect 164923 79792 165108 79794
rect 164923 79736 164928 79792
rect 164984 79736 165108 79792
rect 164923 79734 165108 79736
rect 164804 79732 164810 79734
rect 164693 79731 164759 79732
rect 164923 79731 164989 79734
rect 165102 79732 165108 79734
rect 165172 79794 165178 79796
rect 165172 79734 165584 79794
rect 165172 79732 165178 79734
rect 165524 79661 165584 79734
rect 162158 79658 162164 79660
rect 160940 79656 161032 79658
rect 160982 79600 161032 79656
rect 160940 79598 161032 79600
rect 161844 79598 162164 79658
rect 160940 79596 160987 79598
rect 162158 79596 162164 79598
rect 162228 79596 162234 79660
rect 162442 79656 162551 79661
rect 162442 79600 162490 79656
rect 162546 79600 162551 79656
rect 162442 79598 162551 79600
rect 162718 79656 162827 79661
rect 162718 79600 162766 79656
rect 162822 79600 162827 79656
rect 162718 79598 162827 79600
rect 160921 79595 160987 79596
rect 162485 79595 162551 79598
rect 162761 79595 162827 79598
rect 163078 79596 163084 79660
rect 163148 79658 163154 79660
rect 163221 79658 163287 79661
rect 163148 79656 163287 79658
rect 163148 79600 163226 79656
rect 163282 79600 163287 79656
rect 163148 79598 163287 79600
rect 163148 79596 163154 79598
rect 163221 79595 163287 79598
rect 163630 79596 163636 79660
rect 163700 79658 163706 79660
rect 163773 79658 163839 79661
rect 164233 79660 164299 79661
rect 163700 79656 163839 79658
rect 163700 79600 163778 79656
rect 163834 79600 163839 79656
rect 163700 79598 163839 79600
rect 163700 79596 163706 79598
rect 163773 79595 163839 79598
rect 164182 79596 164188 79660
rect 164252 79658 164299 79660
rect 164252 79656 164344 79658
rect 164294 79600 164344 79656
rect 164252 79598 164344 79600
rect 165521 79656 165587 79661
rect 165521 79600 165526 79656
rect 165582 79600 165587 79656
rect 164252 79596 164299 79598
rect 164233 79595 164299 79596
rect 165521 79595 165587 79600
rect 161606 79460 161612 79524
rect 161676 79522 161682 79524
rect 162209 79522 162275 79525
rect 161676 79520 162275 79522
rect 161676 79464 162214 79520
rect 162270 79464 162275 79520
rect 161676 79462 162275 79464
rect 161676 79460 161682 79462
rect 162209 79459 162275 79462
rect 162342 79460 162348 79524
rect 162412 79522 162418 79524
rect 162669 79522 162735 79525
rect 162412 79520 162735 79522
rect 162412 79464 162674 79520
rect 162730 79464 162735 79520
rect 162412 79462 162735 79464
rect 162412 79460 162418 79462
rect 162669 79459 162735 79462
rect 163262 79460 163268 79524
rect 163332 79522 163338 79524
rect 164049 79522 164115 79525
rect 163332 79520 164115 79522
rect 163332 79464 164054 79520
rect 164110 79464 164115 79520
rect 163332 79462 164115 79464
rect 163332 79460 163338 79462
rect 164049 79459 164115 79462
rect 164550 79460 164556 79524
rect 164620 79522 164626 79524
rect 164785 79522 164851 79525
rect 164620 79520 164851 79522
rect 164620 79464 164790 79520
rect 164846 79464 164851 79520
rect 164620 79462 164851 79464
rect 165662 79522 165722 79901
rect 166027 79872 166032 79928
rect 166088 79872 166093 79928
rect 166027 79867 166093 79872
rect 166488 79870 166580 79930
rect 166574 79868 166580 79870
rect 166644 79868 166650 79932
rect 166942 79930 166948 79932
rect 166856 79870 166948 79930
rect 166942 79868 166948 79870
rect 167012 79868 167018 79932
rect 167131 79930 167197 79933
rect 167088 79928 167197 79930
rect 167088 79872 167136 79928
rect 167192 79872 167197 79928
rect 167499 79928 167565 79933
rect 166579 79867 166645 79868
rect 166947 79867 167013 79868
rect 167088 79867 167197 79872
rect 167315 79894 167381 79899
rect 165889 79794 165955 79797
rect 166022 79794 166028 79796
rect 165889 79792 166028 79794
rect 165889 79736 165894 79792
rect 165950 79736 166028 79792
rect 165889 79734 166028 79736
rect 165889 79731 165955 79734
rect 166022 79732 166028 79734
rect 166092 79732 166098 79796
rect 167088 79661 167148 79867
rect 167315 79838 167320 79894
rect 167376 79838 167381 79894
rect 167499 79872 167504 79928
rect 167560 79872 167565 79928
rect 167499 79867 167565 79872
rect 167732 79906 167780 79962
rect 167836 79906 167841 79962
rect 168235 79964 168301 79967
rect 168235 79962 168358 79964
rect 168051 79932 168117 79933
rect 168235 79932 168240 79962
rect 168296 79932 168358 79962
rect 168046 79930 168052 79932
rect 167732 79901 167841 79906
rect 167315 79833 167381 79838
rect 167318 79661 167378 79833
rect 167502 79796 167562 79867
rect 167494 79732 167500 79796
rect 167564 79732 167570 79796
rect 165838 79596 165844 79660
rect 165908 79658 165914 79660
rect 166625 79658 166691 79661
rect 165908 79656 166691 79658
rect 165908 79600 166630 79656
rect 166686 79600 166691 79656
rect 165908 79598 166691 79600
rect 165908 79596 165914 79598
rect 166625 79595 166691 79598
rect 167085 79656 167151 79661
rect 167085 79600 167090 79656
rect 167146 79600 167151 79656
rect 167085 79595 167151 79600
rect 167269 79656 167378 79661
rect 167269 79600 167274 79656
rect 167330 79600 167378 79656
rect 167269 79598 167378 79600
rect 167545 79658 167611 79661
rect 167732 79658 167792 79901
rect 167960 79870 168052 79930
rect 168046 79868 168052 79870
rect 168116 79868 168122 79932
rect 168230 79868 168236 79932
rect 168300 79904 168358 79932
rect 168300 79868 168306 79904
rect 168051 79867 168117 79868
rect 168422 79831 168482 80142
rect 170078 80142 170260 80202
rect 168598 80004 168604 80068
rect 168668 80066 168674 80068
rect 168668 80006 169034 80066
rect 168668 80004 168674 80006
rect 168787 79928 168853 79933
rect 168787 79872 168792 79928
rect 168848 79872 168853 79928
rect 168787 79867 168853 79872
rect 168974 79930 169034 80006
rect 170078 79967 170138 80142
rect 170254 80140 170260 80142
rect 170324 80140 170330 80204
rect 172830 80140 172836 80204
rect 172900 80202 172906 80204
rect 172900 80142 173404 80202
rect 172900 80140 172906 80142
rect 169155 79962 169221 79967
rect 169155 79930 169160 79962
rect 168974 79906 169160 79930
rect 169216 79906 169221 79962
rect 168974 79901 169221 79906
rect 169431 79964 169497 79967
rect 169431 79962 169540 79964
rect 169431 79906 169436 79962
rect 169492 79906 169540 79962
rect 169431 79901 169540 79906
rect 170075 79962 170141 79967
rect 170075 79906 170080 79962
rect 170136 79906 170141 79962
rect 172743 79964 172809 79967
rect 172927 79964 172993 79967
rect 172743 79962 172852 79964
rect 170075 79901 170141 79906
rect 170443 79930 170509 79933
rect 170990 79930 170996 79932
rect 170443 79928 170996 79930
rect 168974 79870 169218 79901
rect 168419 79826 168485 79831
rect 168419 79770 168424 79826
rect 168480 79770 168485 79826
rect 168419 79765 168485 79770
rect 168790 79794 168850 79867
rect 169017 79794 169083 79797
rect 169334 79794 169340 79796
rect 168790 79792 169340 79794
rect 168790 79736 169022 79792
rect 169078 79736 169340 79792
rect 168790 79734 169340 79736
rect 169017 79731 169083 79734
rect 169334 79732 169340 79734
rect 169404 79732 169410 79796
rect 169480 79794 169540 79901
rect 170443 79872 170448 79928
rect 170504 79872 170996 79928
rect 170443 79870 170996 79872
rect 170443 79867 170509 79870
rect 170990 79868 170996 79870
rect 171060 79868 171066 79932
rect 171271 79930 171337 79933
rect 171547 79932 171613 79933
rect 171542 79930 171548 79932
rect 171271 79928 171380 79930
rect 171271 79872 171276 79928
rect 171332 79872 171380 79928
rect 171271 79867 171380 79872
rect 171456 79870 171548 79930
rect 171542 79868 171548 79870
rect 171612 79868 171618 79932
rect 171726 79868 171732 79932
rect 171796 79930 171802 79932
rect 172099 79930 172165 79933
rect 171796 79928 172165 79930
rect 171796 79872 172104 79928
rect 172160 79872 172165 79928
rect 171796 79870 172165 79872
rect 171796 79868 171802 79870
rect 171547 79867 171613 79868
rect 172099 79867 172165 79870
rect 172283 79930 172349 79933
rect 172283 79928 172392 79930
rect 172283 79872 172288 79928
rect 172344 79872 172392 79928
rect 172743 79906 172748 79962
rect 172804 79906 172852 79962
rect 172743 79901 172852 79906
rect 172927 79962 173036 79964
rect 172927 79906 172932 79962
rect 172988 79932 173036 79962
rect 172988 79906 173020 79932
rect 172927 79901 173020 79906
rect 172283 79867 172392 79872
rect 169702 79794 169708 79796
rect 169480 79734 169708 79794
rect 169702 79732 169708 79734
rect 169772 79732 169778 79796
rect 169886 79732 169892 79796
rect 169956 79794 169962 79796
rect 170995 79794 171061 79797
rect 171174 79794 171180 79796
rect 169956 79792 171180 79794
rect 169956 79736 171000 79792
rect 171056 79736 171180 79792
rect 169956 79734 171180 79736
rect 169956 79732 169962 79734
rect 170995 79731 171061 79734
rect 171174 79732 171180 79734
rect 171244 79732 171250 79796
rect 171320 79794 171380 79867
rect 172094 79794 172100 79796
rect 171320 79734 172100 79794
rect 172094 79732 172100 79734
rect 172164 79732 172170 79796
rect 167545 79656 167792 79658
rect 167545 79600 167550 79656
rect 167606 79600 167792 79656
rect 167545 79598 167792 79600
rect 167269 79595 167335 79598
rect 167545 79595 167611 79598
rect 167862 79596 167868 79660
rect 167932 79658 167938 79660
rect 168005 79658 168071 79661
rect 169150 79658 169156 79660
rect 167932 79656 168071 79658
rect 167932 79600 168010 79656
rect 168066 79600 168071 79656
rect 167932 79598 168071 79600
rect 167932 79596 167938 79598
rect 168005 79595 168071 79598
rect 168790 79598 169156 79658
rect 166758 79522 166764 79524
rect 165662 79462 166764 79522
rect 164620 79460 164626 79462
rect 164785 79459 164851 79462
rect 166758 79460 166764 79462
rect 166828 79460 166834 79524
rect 167310 79460 167316 79524
rect 167380 79522 167386 79524
rect 167453 79522 167519 79525
rect 167380 79520 167519 79522
rect 167380 79464 167458 79520
rect 167514 79464 167519 79520
rect 167380 79462 167519 79464
rect 167380 79460 167386 79462
rect 167453 79459 167519 79462
rect 167678 79460 167684 79524
rect 167748 79522 167754 79524
rect 168005 79522 168071 79525
rect 167748 79520 168071 79522
rect 167748 79464 168010 79520
rect 168066 79464 168071 79520
rect 167748 79462 168071 79464
rect 167748 79460 167754 79462
rect 168005 79459 168071 79462
rect 168373 79522 168439 79525
rect 168790 79522 168850 79598
rect 169150 79596 169156 79598
rect 169220 79658 169226 79660
rect 169385 79658 169451 79661
rect 169220 79656 169451 79658
rect 169220 79600 169390 79656
rect 169446 79600 169451 79656
rect 169220 79598 169451 79600
rect 169220 79596 169226 79598
rect 169385 79595 169451 79598
rect 170070 79596 170076 79660
rect 170140 79658 170146 79660
rect 170857 79658 170923 79661
rect 170140 79656 170923 79658
rect 170140 79600 170862 79656
rect 170918 79600 170923 79656
rect 170140 79598 170923 79600
rect 170140 79596 170146 79598
rect 170857 79595 170923 79598
rect 171358 79596 171364 79660
rect 171428 79658 171434 79660
rect 171869 79658 171935 79661
rect 171428 79656 171935 79658
rect 171428 79600 171874 79656
rect 171930 79600 171935 79656
rect 171428 79598 171935 79600
rect 171428 79596 171434 79598
rect 171869 79595 171935 79598
rect 168373 79520 168850 79522
rect 168373 79464 168378 79520
rect 168434 79464 168850 79520
rect 168373 79462 168850 79464
rect 169201 79522 169267 79525
rect 169518 79522 169524 79524
rect 169201 79520 169524 79522
rect 169201 79464 169206 79520
rect 169262 79464 169524 79520
rect 169201 79462 169524 79464
rect 168373 79459 168439 79462
rect 169201 79459 169267 79462
rect 169518 79460 169524 79462
rect 169588 79460 169594 79524
rect 170622 79460 170628 79524
rect 170692 79522 170698 79524
rect 171041 79522 171107 79525
rect 171685 79522 171751 79525
rect 170692 79520 171107 79522
rect 170692 79464 171046 79520
rect 171102 79464 171107 79520
rect 170692 79462 171107 79464
rect 170692 79460 170698 79462
rect 171041 79459 171107 79462
rect 171320 79520 171751 79522
rect 171320 79464 171690 79520
rect 171746 79464 171751 79520
rect 171320 79462 171751 79464
rect 159950 79324 159956 79388
rect 160020 79386 160026 79388
rect 169385 79386 169451 79389
rect 160020 79384 169451 79386
rect 160020 79328 169390 79384
rect 169446 79328 169451 79384
rect 160020 79326 169451 79328
rect 160020 79324 160026 79326
rect 169385 79323 169451 79326
rect 170305 79386 170371 79389
rect 170438 79386 170444 79388
rect 170305 79384 170444 79386
rect 170305 79328 170310 79384
rect 170366 79328 170444 79384
rect 170305 79326 170444 79328
rect 170305 79323 170371 79326
rect 170438 79324 170444 79326
rect 170508 79324 170514 79388
rect 163497 79250 163563 79253
rect 163998 79250 164004 79252
rect 163497 79248 164004 79250
rect 163497 79192 163502 79248
rect 163558 79192 164004 79248
rect 163497 79190 164004 79192
rect 163497 79187 163563 79190
rect 163998 79188 164004 79190
rect 164068 79188 164074 79252
rect 164918 79188 164924 79252
rect 164988 79250 164994 79252
rect 165245 79250 165311 79253
rect 164988 79248 165311 79250
rect 164988 79192 165250 79248
rect 165306 79192 165311 79248
rect 164988 79190 165311 79192
rect 164988 79188 164994 79190
rect 165245 79187 165311 79190
rect 166206 79188 166212 79252
rect 166276 79250 166282 79252
rect 166993 79250 167059 79253
rect 166276 79248 167059 79250
rect 166276 79192 166998 79248
rect 167054 79192 167059 79248
rect 166276 79190 167059 79192
rect 166276 79188 166282 79190
rect 166993 79187 167059 79190
rect 169017 79250 169083 79253
rect 171320 79250 171380 79462
rect 171685 79459 171751 79462
rect 172053 79522 172119 79525
rect 172332 79522 172392 79867
rect 172792 79794 172852 79901
rect 172976 79870 173020 79901
rect 173014 79868 173020 79870
rect 173084 79868 173090 79932
rect 173344 79930 173404 80142
rect 175590 80140 175596 80204
rect 175660 80202 175666 80204
rect 175660 80142 176210 80202
rect 175660 80140 175666 80142
rect 176150 80066 176210 80142
rect 176326 80140 176332 80204
rect 176396 80202 176402 80204
rect 181437 80202 181503 80205
rect 176396 80200 181503 80202
rect 176396 80144 181442 80200
rect 181498 80144 181503 80200
rect 176396 80142 181503 80144
rect 186270 80202 186330 80278
rect 186865 80202 186931 80205
rect 187417 80202 187483 80205
rect 186270 80200 187483 80202
rect 186270 80144 186870 80200
rect 186926 80144 187422 80200
rect 187478 80144 187483 80200
rect 186270 80142 187483 80144
rect 176396 80140 176402 80142
rect 181437 80139 181503 80142
rect 186865 80139 186931 80142
rect 187417 80139 187483 80142
rect 179321 80066 179387 80069
rect 186262 80066 186268 80068
rect 176150 80006 176716 80066
rect 173847 79962 173913 79967
rect 173479 79930 173545 79933
rect 173344 79928 173545 79930
rect 173344 79872 173484 79928
rect 173540 79872 173545 79928
rect 173847 79906 173852 79962
rect 173908 79906 173913 79962
rect 173847 79901 173913 79906
rect 174307 79930 174373 79933
rect 174854 79930 174860 79932
rect 174307 79928 174860 79930
rect 173344 79870 173545 79872
rect 173479 79867 173545 79870
rect 173014 79794 173020 79796
rect 172792 79734 173020 79794
rect 173014 79732 173020 79734
rect 173084 79732 173090 79796
rect 173566 79732 173572 79796
rect 173636 79794 173642 79796
rect 173850 79794 173910 79901
rect 174307 79872 174312 79928
rect 174368 79872 174860 79928
rect 174307 79870 174860 79872
rect 174307 79867 174373 79870
rect 174854 79868 174860 79870
rect 174924 79868 174930 79932
rect 175038 79868 175044 79932
rect 175108 79930 175114 79932
rect 175227 79930 175293 79933
rect 175411 79930 175477 79933
rect 175108 79928 175293 79930
rect 175108 79872 175232 79928
rect 175288 79872 175293 79928
rect 175108 79870 175293 79872
rect 175108 79868 175114 79870
rect 175227 79867 175293 79870
rect 175368 79928 175477 79930
rect 175368 79872 175416 79928
rect 175472 79872 175477 79928
rect 175368 79867 175477 79872
rect 175590 79868 175596 79932
rect 175660 79930 175666 79932
rect 175779 79930 175845 79933
rect 176331 79932 176397 79933
rect 175660 79928 175845 79930
rect 175660 79872 175784 79928
rect 175840 79872 175845 79928
rect 175660 79870 175845 79872
rect 175660 79868 175666 79870
rect 175779 79867 175845 79870
rect 176142 79868 176148 79932
rect 176212 79930 176218 79932
rect 176212 79868 176256 79930
rect 176326 79868 176332 79932
rect 176396 79930 176402 79932
rect 176396 79870 176488 79930
rect 176396 79868 176402 79870
rect 173636 79734 173910 79794
rect 173636 79732 173642 79734
rect 174118 79732 174124 79796
rect 174188 79794 174194 79796
rect 174537 79794 174603 79797
rect 174188 79792 174603 79794
rect 174188 79736 174542 79792
rect 174598 79736 174603 79792
rect 174188 79734 174603 79736
rect 174188 79732 174194 79734
rect 174537 79731 174603 79734
rect 174670 79732 174676 79796
rect 174740 79794 174746 79796
rect 175135 79794 175201 79797
rect 174740 79792 175201 79794
rect 174740 79736 175140 79792
rect 175196 79736 175201 79792
rect 174740 79734 175201 79736
rect 175368 79794 175428 79867
rect 176196 79797 176256 79868
rect 176331 79867 176397 79868
rect 175958 79794 175964 79796
rect 175368 79734 175964 79794
rect 174740 79732 174746 79734
rect 175135 79731 175201 79734
rect 175958 79732 175964 79734
rect 176028 79732 176034 79796
rect 176193 79792 176259 79797
rect 176193 79736 176198 79792
rect 176254 79736 176259 79792
rect 176193 79731 176259 79736
rect 176515 79794 176581 79797
rect 176656 79794 176716 80006
rect 179321 80064 186268 80066
rect 179321 80008 179326 80064
rect 179382 80008 186268 80064
rect 179321 80006 186268 80008
rect 179321 80003 179387 80006
rect 186262 80004 186268 80006
rect 186332 80004 186338 80068
rect 177343 79964 177409 79967
rect 177300 79962 177409 79964
rect 177062 79868 177068 79932
rect 177132 79930 177138 79932
rect 177300 79930 177348 79962
rect 177132 79906 177348 79930
rect 177404 79906 177409 79962
rect 177132 79901 177409 79906
rect 177527 79964 177593 79967
rect 177527 79962 177636 79964
rect 177527 79906 177532 79962
rect 177588 79932 177636 79962
rect 177588 79906 177620 79932
rect 177527 79901 177620 79906
rect 177132 79870 177360 79901
rect 177576 79870 177620 79901
rect 177132 79868 177138 79870
rect 177614 79868 177620 79870
rect 177684 79868 177690 79932
rect 176515 79792 176716 79794
rect 176515 79736 176520 79792
rect 176576 79736 176716 79792
rect 176515 79734 176716 79736
rect 176515 79731 176581 79734
rect 176878 79732 176884 79796
rect 176948 79794 176954 79796
rect 177481 79794 177547 79797
rect 182081 79794 182147 79797
rect 176948 79792 182147 79794
rect 176948 79736 177486 79792
rect 177542 79736 182086 79792
rect 182142 79736 182147 79792
rect 176948 79734 182147 79736
rect 176948 79732 176954 79734
rect 177481 79731 177547 79734
rect 182081 79731 182147 79734
rect 173249 79658 173315 79661
rect 173382 79658 173388 79660
rect 173249 79656 173388 79658
rect 173249 79600 173254 79656
rect 173310 79600 173388 79656
rect 173249 79598 173388 79600
rect 173249 79595 173315 79598
rect 173382 79596 173388 79598
rect 173452 79596 173458 79660
rect 174302 79596 174308 79660
rect 174372 79658 174378 79660
rect 174813 79658 174879 79661
rect 174372 79656 174879 79658
rect 174372 79600 174818 79656
rect 174874 79600 174879 79656
rect 174372 79598 174879 79600
rect 174372 79596 174378 79598
rect 174813 79595 174879 79598
rect 175273 79658 175339 79661
rect 175774 79658 175780 79660
rect 175273 79656 175780 79658
rect 175273 79600 175278 79656
rect 175334 79600 175780 79656
rect 175273 79598 175780 79600
rect 175273 79595 175339 79598
rect 175774 79596 175780 79598
rect 175844 79596 175850 79660
rect 176101 79658 176167 79661
rect 176101 79656 186330 79658
rect 176101 79600 176106 79656
rect 176162 79600 186330 79656
rect 176101 79598 186330 79600
rect 176101 79595 176167 79598
rect 172053 79520 172392 79522
rect 172053 79464 172058 79520
rect 172114 79464 172392 79520
rect 172053 79462 172392 79464
rect 172053 79459 172119 79462
rect 172646 79460 172652 79524
rect 172716 79522 172722 79524
rect 173249 79522 173315 79525
rect 173709 79522 173775 79525
rect 172716 79520 173775 79522
rect 172716 79464 173254 79520
rect 173310 79464 173714 79520
rect 173770 79464 173775 79520
rect 172716 79462 173775 79464
rect 172716 79460 172722 79462
rect 173249 79459 173315 79462
rect 173709 79459 173775 79462
rect 174077 79522 174143 79525
rect 175181 79522 175247 79525
rect 174077 79520 175247 79522
rect 174077 79464 174082 79520
rect 174138 79464 175186 79520
rect 175242 79464 175247 79520
rect 174077 79462 175247 79464
rect 174077 79459 174143 79462
rect 175181 79459 175247 79462
rect 175406 79460 175412 79524
rect 175476 79522 175482 79524
rect 175917 79522 175983 79525
rect 175476 79520 175983 79522
rect 175476 79464 175922 79520
rect 175978 79464 175983 79520
rect 175476 79462 175983 79464
rect 175476 79460 175482 79462
rect 175917 79459 175983 79462
rect 176653 79522 176719 79525
rect 177062 79522 177068 79524
rect 176653 79520 177068 79522
rect 176653 79464 176658 79520
rect 176714 79464 177068 79520
rect 176653 79462 177068 79464
rect 176653 79459 176719 79462
rect 177062 79460 177068 79462
rect 177132 79460 177138 79524
rect 177665 79522 177731 79525
rect 177798 79522 177804 79524
rect 177665 79520 177804 79522
rect 177665 79464 177670 79520
rect 177726 79464 177804 79520
rect 177665 79462 177804 79464
rect 177665 79459 177731 79462
rect 177798 79460 177804 79462
rect 177868 79460 177874 79524
rect 180926 79460 180932 79524
rect 180996 79522 181002 79524
rect 181069 79522 181135 79525
rect 180996 79520 181135 79522
rect 180996 79464 181074 79520
rect 181130 79464 181135 79520
rect 180996 79462 181135 79464
rect 180996 79460 181002 79462
rect 181069 79459 181135 79462
rect 186270 79386 186330 79598
rect 193990 79386 193996 79388
rect 171688 79326 183570 79386
rect 186270 79326 193996 79386
rect 171688 79253 171748 79326
rect 169017 79248 171380 79250
rect 169017 79192 169022 79248
rect 169078 79192 171380 79248
rect 169017 79190 171380 79192
rect 171501 79250 171567 79253
rect 171685 79250 171751 79253
rect 171501 79248 171751 79250
rect 171501 79192 171506 79248
rect 171562 79192 171690 79248
rect 171746 79192 171751 79248
rect 171501 79190 171751 79192
rect 169017 79187 169083 79190
rect 171501 79187 171567 79190
rect 171685 79187 171751 79190
rect 171910 79188 171916 79252
rect 171980 79250 171986 79252
rect 172329 79250 172395 79253
rect 171980 79248 172395 79250
rect 171980 79192 172334 79248
rect 172390 79192 172395 79248
rect 171980 79190 172395 79192
rect 171980 79188 171986 79190
rect 172329 79187 172395 79190
rect 173065 79250 173131 79253
rect 175222 79250 175228 79252
rect 173065 79248 175228 79250
rect 173065 79192 173070 79248
rect 173126 79192 175228 79248
rect 173065 79190 175228 79192
rect 173065 79187 173131 79190
rect 175222 79188 175228 79190
rect 175292 79188 175298 79252
rect 175958 79188 175964 79252
rect 176028 79250 176034 79252
rect 177573 79250 177639 79253
rect 176028 79248 177639 79250
rect 176028 79192 177578 79248
rect 177634 79192 177639 79248
rect 176028 79190 177639 79192
rect 183510 79250 183570 79326
rect 193990 79324 193996 79326
rect 194060 79324 194066 79388
rect 190862 79250 190868 79252
rect 183510 79190 190868 79250
rect 176028 79188 176034 79190
rect 177573 79187 177639 79190
rect 190862 79188 190868 79190
rect 190932 79188 190938 79252
rect 160185 79114 160251 79117
rect 150084 79112 160251 79114
rect 150084 79056 160190 79112
rect 160246 79056 160251 79112
rect 150084 79054 160251 79056
rect 150084 79052 150090 79054
rect 160185 79051 160251 79054
rect 160553 79114 160619 79117
rect 160686 79114 160692 79116
rect 160553 79112 160692 79114
rect 160553 79056 160558 79112
rect 160614 79056 160692 79112
rect 160553 79054 160692 79056
rect 160553 79051 160619 79054
rect 160686 79052 160692 79054
rect 160756 79052 160762 79116
rect 161841 79114 161907 79117
rect 162526 79114 162532 79116
rect 161841 79112 162532 79114
rect 161841 79056 161846 79112
rect 161902 79056 162532 79112
rect 161841 79054 162532 79056
rect 161841 79051 161907 79054
rect 162526 79052 162532 79054
rect 162596 79052 162602 79116
rect 165705 79114 165771 79117
rect 166942 79114 166948 79116
rect 165705 79112 166948 79114
rect 165705 79056 165710 79112
rect 165766 79056 166948 79112
rect 165705 79054 166948 79056
rect 165705 79051 165771 79054
rect 166942 79052 166948 79054
rect 167012 79114 167018 79116
rect 167361 79114 167427 79117
rect 167012 79112 167427 79114
rect 167012 79056 167366 79112
rect 167422 79056 167427 79112
rect 167012 79054 167427 79056
rect 167012 79052 167018 79054
rect 167361 79051 167427 79054
rect 167545 79114 167611 79117
rect 167862 79114 167868 79116
rect 167545 79112 167868 79114
rect 167545 79056 167550 79112
rect 167606 79056 167868 79112
rect 167545 79054 167868 79056
rect 167545 79051 167611 79054
rect 167862 79052 167868 79054
rect 167932 79052 167938 79116
rect 168966 79052 168972 79116
rect 169036 79114 169042 79116
rect 169753 79114 169819 79117
rect 169036 79112 169819 79114
rect 169036 79056 169758 79112
rect 169814 79056 169819 79112
rect 169036 79054 169819 79056
rect 169036 79052 169042 79054
rect 169753 79051 169819 79054
rect 170489 79114 170555 79117
rect 170806 79114 170812 79116
rect 170489 79112 170812 79114
rect 170489 79056 170494 79112
rect 170550 79056 170812 79112
rect 170489 79054 170812 79056
rect 170489 79051 170555 79054
rect 170806 79052 170812 79054
rect 170876 79052 170882 79116
rect 173198 79114 173204 79116
rect 171964 79054 173204 79114
rect 125244 78918 139410 78978
rect 139577 78978 139643 78981
rect 140446 78978 140452 78980
rect 139577 78976 140452 78978
rect 139577 78920 139582 78976
rect 139638 78920 140452 78976
rect 139577 78918 140452 78920
rect 125244 78916 125250 78918
rect 139577 78915 139643 78918
rect 140446 78916 140452 78918
rect 140516 78978 140522 78980
rect 140681 78978 140747 78981
rect 140516 78976 140747 78978
rect 140516 78920 140686 78976
rect 140742 78920 140747 78976
rect 140516 78918 140747 78920
rect 140516 78916 140522 78918
rect 140681 78915 140747 78918
rect 140865 78978 140931 78981
rect 142102 78978 142108 78980
rect 140865 78976 142108 78978
rect 140865 78920 140870 78976
rect 140926 78920 142108 78976
rect 140865 78918 142108 78920
rect 140865 78915 140931 78918
rect 142102 78916 142108 78918
rect 142172 78978 142178 78980
rect 142654 78978 142660 78980
rect 142172 78918 142660 78978
rect 142172 78916 142178 78918
rect 142654 78916 142660 78918
rect 142724 78916 142730 78980
rect 143206 78916 143212 78980
rect 143276 78978 143282 78980
rect 143809 78978 143875 78981
rect 143276 78976 143875 78978
rect 143276 78920 143814 78976
rect 143870 78920 143875 78976
rect 143276 78918 143875 78920
rect 143276 78916 143282 78918
rect 143809 78915 143875 78918
rect 145598 78916 145604 78980
rect 145668 78978 145674 78980
rect 161841 78978 161907 78981
rect 145668 78976 161907 78978
rect 145668 78920 161846 78976
rect 161902 78920 161907 78976
rect 145668 78918 161907 78920
rect 145668 78916 145674 78918
rect 161841 78915 161907 78918
rect 170489 78978 170555 78981
rect 170990 78978 170996 78980
rect 170489 78976 170996 78978
rect 170489 78920 170494 78976
rect 170550 78920 170996 78976
rect 170489 78918 170996 78920
rect 170489 78915 170555 78918
rect 170990 78916 170996 78918
rect 171060 78916 171066 78980
rect 171225 78978 171291 78981
rect 171964 78978 172024 79054
rect 173198 79052 173204 79054
rect 173268 79052 173274 79116
rect 173341 79114 173407 79117
rect 195053 79114 195119 79117
rect 173341 79112 195119 79114
rect 173341 79056 173346 79112
rect 173402 79056 195058 79112
rect 195114 79056 195119 79112
rect 173341 79054 195119 79056
rect 173341 79051 173407 79054
rect 195053 79051 195119 79054
rect 171225 78976 172024 78978
rect 171225 78920 171230 78976
rect 171286 78920 172024 78976
rect 171225 78918 172024 78920
rect 171225 78915 171291 78918
rect 172094 78916 172100 78980
rect 172164 78978 172170 78980
rect 172237 78978 172303 78981
rect 172164 78976 172303 78978
rect 172164 78920 172242 78976
rect 172298 78920 172303 78976
rect 172164 78918 172303 78920
rect 172164 78916 172170 78918
rect 172237 78915 172303 78918
rect 175733 78978 175799 78981
rect 179505 78980 179571 78981
rect 176510 78978 176516 78980
rect 175733 78976 176516 78978
rect 175733 78920 175738 78976
rect 175794 78920 176516 78976
rect 175733 78918 176516 78920
rect 175733 78915 175799 78918
rect 176510 78916 176516 78918
rect 176580 78916 176586 78980
rect 179454 78978 179460 78980
rect 179414 78918 179460 78978
rect 179524 78976 179571 78980
rect 179566 78920 179571 78976
rect 179454 78916 179460 78918
rect 179524 78916 179571 78920
rect 180742 78916 180748 78980
rect 180812 78978 180818 78980
rect 180885 78978 180951 78981
rect 180812 78976 180951 78978
rect 180812 78920 180890 78976
rect 180946 78920 180951 78976
rect 180812 78918 180951 78920
rect 180812 78916 180818 78918
rect 179505 78915 179571 78916
rect 180885 78915 180951 78918
rect 181161 78978 181227 78981
rect 197997 78978 198063 78981
rect 181161 78976 198063 78978
rect 181161 78920 181166 78976
rect 181222 78920 198002 78976
rect 198058 78920 198063 78976
rect 181161 78918 198063 78920
rect 181161 78915 181227 78918
rect 197997 78915 198063 78918
rect 198958 78916 198964 78980
rect 199028 78978 199034 78980
rect 199326 78978 199332 78980
rect 199028 78918 199332 78978
rect 199028 78916 199034 78918
rect 199326 78916 199332 78918
rect 199396 78978 199402 78980
rect 536833 78978 536899 78981
rect 199396 78976 536899 78978
rect 199396 78920 536838 78976
rect 536894 78920 536899 78976
rect 199396 78918 536899 78920
rect 199396 78916 199402 78918
rect 536833 78915 536899 78918
rect 124070 78780 124076 78844
rect 124140 78842 124146 78844
rect 124140 78782 147690 78842
rect 124140 78780 124146 78782
rect 130878 78644 130884 78708
rect 130948 78706 130954 78708
rect 138289 78706 138355 78709
rect 130948 78704 138355 78706
rect 130948 78648 138294 78704
rect 138350 78648 138355 78704
rect 130948 78646 138355 78648
rect 130948 78644 130954 78646
rect 138289 78643 138355 78646
rect 138614 78646 139226 78706
rect 124806 78508 124812 78572
rect 124876 78570 124882 78572
rect 130837 78570 130903 78573
rect 132861 78572 132927 78573
rect 132861 78570 132908 78572
rect 124876 78568 130903 78570
rect 124876 78512 130842 78568
rect 130898 78512 130903 78568
rect 124876 78510 130903 78512
rect 132816 78568 132908 78570
rect 132816 78512 132866 78568
rect 132816 78510 132908 78512
rect 124876 78508 124882 78510
rect 130837 78507 130903 78510
rect 132861 78508 132908 78510
rect 132972 78508 132978 78572
rect 133045 78570 133111 78573
rect 133454 78570 133460 78572
rect 133045 78568 133460 78570
rect 133045 78512 133050 78568
rect 133106 78512 133460 78568
rect 133045 78510 133460 78512
rect 132861 78507 132927 78508
rect 133045 78507 133111 78510
rect 133454 78508 133460 78510
rect 133524 78508 133530 78572
rect 135621 78570 135687 78573
rect 135846 78570 135852 78572
rect 135621 78568 135852 78570
rect 135621 78512 135626 78568
rect 135682 78512 135852 78568
rect 135621 78510 135852 78512
rect 135621 78507 135687 78510
rect 135846 78508 135852 78510
rect 135916 78508 135922 78572
rect 137134 78508 137140 78572
rect 137204 78570 137210 78572
rect 137921 78570 137987 78573
rect 138105 78572 138171 78573
rect 137204 78568 137987 78570
rect 137204 78512 137926 78568
rect 137982 78512 137987 78568
rect 137204 78510 137987 78512
rect 137204 78508 137210 78510
rect 137921 78507 137987 78510
rect 138054 78508 138060 78572
rect 138124 78570 138171 78572
rect 138614 78570 138674 78646
rect 138124 78568 138216 78570
rect 138166 78512 138216 78568
rect 138124 78510 138216 78512
rect 138430 78510 138674 78570
rect 139166 78570 139226 78646
rect 139342 78644 139348 78708
rect 139412 78706 139418 78708
rect 139669 78706 139735 78709
rect 139412 78704 139735 78706
rect 139412 78648 139674 78704
rect 139730 78648 139735 78704
rect 139412 78646 139735 78648
rect 139412 78644 139418 78646
rect 139669 78643 139735 78646
rect 143390 78644 143396 78708
rect 143460 78706 143466 78708
rect 143717 78706 143783 78709
rect 143460 78704 143783 78706
rect 143460 78648 143722 78704
rect 143778 78648 143783 78704
rect 143460 78646 143783 78648
rect 147630 78706 147690 78782
rect 148910 78780 148916 78844
rect 148980 78842 148986 78844
rect 161657 78842 161723 78845
rect 148980 78840 161723 78842
rect 148980 78784 161662 78840
rect 161718 78784 161723 78840
rect 148980 78782 161723 78784
rect 148980 78780 148986 78782
rect 161657 78779 161723 78782
rect 162209 78842 162275 78845
rect 382273 78842 382339 78845
rect 162209 78840 382339 78842
rect 162209 78784 162214 78840
rect 162270 78784 382278 78840
rect 382334 78784 382339 78840
rect 162209 78782 382339 78784
rect 162209 78779 162275 78782
rect 382273 78779 382339 78782
rect 151169 78706 151235 78709
rect 151486 78706 151492 78708
rect 147630 78646 150634 78706
rect 143460 78644 143466 78646
rect 143717 78643 143783 78646
rect 146753 78570 146819 78573
rect 139166 78568 146819 78570
rect 139166 78512 146758 78568
rect 146814 78512 146819 78568
rect 139166 78510 146819 78512
rect 150574 78570 150634 78646
rect 151169 78704 151492 78706
rect 151169 78648 151174 78704
rect 151230 78648 151492 78704
rect 151169 78646 151492 78648
rect 151169 78643 151235 78646
rect 151486 78644 151492 78646
rect 151556 78644 151562 78708
rect 156965 78706 157031 78709
rect 158161 78708 158227 78709
rect 158529 78708 158595 78709
rect 151862 78704 157031 78706
rect 151862 78648 156970 78704
rect 157026 78648 157031 78704
rect 151862 78646 157031 78648
rect 151862 78570 151922 78646
rect 156965 78643 157031 78646
rect 158110 78644 158116 78708
rect 158180 78706 158227 78708
rect 158478 78706 158484 78708
rect 158180 78704 158272 78706
rect 158222 78648 158272 78704
rect 158180 78646 158272 78648
rect 158438 78646 158484 78706
rect 158548 78704 158595 78708
rect 158590 78648 158595 78704
rect 158180 78644 158227 78646
rect 158478 78644 158484 78646
rect 158548 78644 158595 78648
rect 159582 78644 159588 78708
rect 159652 78706 159658 78708
rect 160461 78706 160527 78709
rect 168281 78708 168347 78709
rect 168230 78706 168236 78708
rect 159652 78704 160527 78706
rect 159652 78648 160466 78704
rect 160522 78648 160527 78704
rect 159652 78646 160527 78648
rect 168190 78646 168236 78706
rect 168300 78704 168347 78708
rect 436093 78706 436159 78709
rect 168342 78648 168347 78704
rect 159652 78644 159658 78646
rect 158161 78643 158227 78644
rect 158529 78643 158595 78644
rect 160461 78643 160527 78646
rect 168230 78644 168236 78646
rect 168300 78644 168347 78648
rect 168281 78643 168347 78644
rect 168422 78704 436159 78706
rect 168422 78648 436098 78704
rect 436154 78648 436159 78704
rect 168422 78646 436159 78648
rect 152365 78572 152431 78573
rect 154021 78572 154087 78573
rect 154481 78572 154547 78573
rect 152365 78570 152412 78572
rect 150574 78510 151922 78570
rect 152320 78568 152412 78570
rect 152320 78512 152370 78568
rect 152320 78510 152412 78512
rect 138124 78508 138171 78510
rect 138105 78507 138171 78508
rect 128118 78372 128124 78436
rect 128188 78434 128194 78436
rect 132953 78434 133019 78437
rect 138430 78434 138490 78510
rect 146753 78507 146819 78510
rect 152365 78508 152412 78510
rect 152476 78508 152482 78572
rect 154021 78568 154068 78572
rect 154132 78570 154138 78572
rect 154430 78570 154436 78572
rect 154021 78512 154026 78568
rect 154021 78508 154068 78512
rect 154132 78510 154178 78570
rect 154390 78510 154436 78570
rect 154500 78568 154547 78572
rect 154542 78512 154547 78568
rect 154132 78508 154138 78510
rect 154430 78508 154436 78510
rect 154500 78508 154547 78512
rect 152365 78507 152431 78508
rect 154021 78507 154087 78508
rect 154481 78507 154547 78508
rect 155125 78570 155191 78573
rect 155718 78570 155724 78572
rect 155125 78568 155724 78570
rect 155125 78512 155130 78568
rect 155186 78512 155724 78568
rect 155125 78510 155724 78512
rect 155125 78507 155191 78510
rect 155718 78508 155724 78510
rect 155788 78508 155794 78572
rect 166625 78570 166691 78573
rect 168422 78570 168482 78646
rect 436093 78643 436159 78646
rect 166625 78568 168482 78570
rect 166625 78512 166630 78568
rect 166686 78512 168482 78568
rect 166625 78510 168482 78512
rect 166625 78507 166691 78510
rect 171910 78508 171916 78572
rect 171980 78570 171986 78572
rect 172421 78570 172487 78573
rect 171980 78568 172487 78570
rect 171980 78512 172426 78568
rect 172482 78512 172487 78568
rect 171980 78510 172487 78512
rect 171980 78508 171986 78510
rect 172421 78507 172487 78510
rect 173382 78508 173388 78572
rect 173452 78570 173458 78572
rect 173709 78570 173775 78573
rect 174813 78572 174879 78573
rect 174813 78570 174860 78572
rect 173452 78568 173775 78570
rect 173452 78512 173714 78568
rect 173770 78512 173775 78568
rect 173452 78510 173775 78512
rect 174768 78568 174860 78570
rect 174768 78512 174818 78568
rect 174768 78510 174860 78512
rect 173452 78508 173458 78510
rect 173709 78507 173775 78510
rect 174813 78508 174860 78510
rect 174924 78508 174930 78572
rect 177614 78508 177620 78572
rect 177684 78570 177690 78572
rect 580993 78570 581059 78573
rect 177684 78568 581059 78570
rect 177684 78512 580998 78568
rect 581054 78512 581059 78568
rect 177684 78510 581059 78512
rect 177684 78508 177690 78510
rect 174813 78507 174879 78508
rect 580993 78507 581059 78510
rect 142470 78434 142476 78436
rect 128188 78432 133019 78434
rect 128188 78376 132958 78432
rect 133014 78376 133019 78432
rect 128188 78374 133019 78376
rect 128188 78372 128194 78374
rect 132953 78371 133019 78374
rect 133094 78374 138490 78434
rect 139166 78374 142476 78434
rect 126830 78236 126836 78300
rect 126900 78298 126906 78300
rect 133094 78298 133154 78374
rect 126900 78238 133154 78298
rect 126900 78236 126906 78238
rect 135478 78236 135484 78300
rect 135548 78298 135554 78300
rect 135989 78298 136055 78301
rect 135548 78296 136055 78298
rect 135548 78240 135994 78296
rect 136050 78240 136055 78296
rect 135548 78238 136055 78240
rect 135548 78236 135554 78238
rect 135989 78235 136055 78238
rect 137277 78298 137343 78301
rect 139166 78298 139226 78374
rect 142470 78372 142476 78374
rect 142540 78372 142546 78436
rect 150750 78372 150756 78436
rect 150820 78434 150826 78436
rect 151721 78434 151787 78437
rect 150820 78432 151787 78434
rect 150820 78376 151726 78432
rect 151782 78376 151787 78432
rect 150820 78374 151787 78376
rect 150820 78372 150826 78374
rect 151721 78371 151787 78374
rect 156638 78372 156644 78436
rect 156708 78434 156714 78436
rect 156781 78434 156847 78437
rect 156708 78432 156847 78434
rect 156708 78376 156786 78432
rect 156842 78376 156847 78432
rect 156708 78374 156847 78376
rect 156708 78372 156714 78374
rect 156781 78371 156847 78374
rect 159030 78372 159036 78436
rect 159100 78434 159106 78436
rect 160001 78434 160067 78437
rect 159100 78432 160067 78434
rect 159100 78376 160006 78432
rect 160062 78376 160067 78432
rect 159100 78374 160067 78376
rect 159100 78372 159106 78374
rect 160001 78371 160067 78374
rect 173014 78372 173020 78436
rect 173084 78434 173090 78436
rect 187918 78434 187924 78436
rect 173084 78374 187924 78434
rect 173084 78372 173090 78374
rect 187918 78372 187924 78374
rect 187988 78372 187994 78436
rect 137277 78296 139226 78298
rect 137277 78240 137282 78296
rect 137338 78240 139226 78296
rect 137277 78238 139226 78240
rect 137277 78235 137343 78238
rect 148358 78236 148364 78300
rect 148428 78298 148434 78300
rect 148777 78298 148843 78301
rect 148428 78296 148843 78298
rect 148428 78240 148782 78296
rect 148838 78240 148843 78296
rect 148428 78238 148843 78240
rect 148428 78236 148434 78238
rect 148777 78235 148843 78238
rect 149094 78236 149100 78300
rect 149164 78298 149170 78300
rect 150157 78298 150223 78301
rect 149164 78296 150223 78298
rect 149164 78240 150162 78296
rect 150218 78240 150223 78296
rect 149164 78238 150223 78240
rect 149164 78236 149170 78238
rect 150157 78235 150223 78238
rect 152406 78236 152412 78300
rect 152476 78298 152482 78300
rect 153009 78298 153075 78301
rect 152476 78296 153075 78298
rect 152476 78240 153014 78296
rect 153070 78240 153075 78296
rect 152476 78238 153075 78240
rect 152476 78236 152482 78238
rect 153009 78235 153075 78238
rect 168598 78236 168604 78300
rect 168668 78298 168674 78300
rect 168925 78298 168991 78301
rect 168668 78296 168991 78298
rect 168668 78240 168930 78296
rect 168986 78240 168991 78296
rect 168668 78238 168991 78240
rect 168668 78236 168674 78238
rect 168925 78235 168991 78238
rect 171542 78236 171548 78300
rect 171612 78298 171618 78300
rect 171869 78298 171935 78301
rect 171612 78296 171935 78298
rect 171612 78240 171874 78296
rect 171930 78240 171935 78296
rect 171612 78238 171935 78240
rect 171612 78236 171618 78238
rect 171869 78235 171935 78238
rect 175181 78298 175247 78301
rect 175181 78296 176210 78298
rect 175181 78240 175186 78296
rect 175242 78240 176210 78296
rect 175181 78238 176210 78240
rect 175181 78235 175247 78238
rect 130009 78162 130075 78165
rect 132585 78162 132651 78165
rect 130009 78160 132651 78162
rect 130009 78104 130014 78160
rect 130070 78104 132590 78160
rect 132646 78104 132651 78160
rect 130009 78102 132651 78104
rect 130009 78099 130075 78102
rect 132585 78099 132651 78102
rect 132953 78162 133019 78165
rect 139301 78162 139367 78165
rect 150065 78162 150131 78165
rect 132953 78160 139367 78162
rect 132953 78104 132958 78160
rect 133014 78104 139306 78160
rect 139362 78104 139367 78160
rect 132953 78102 139367 78104
rect 132953 78099 133019 78102
rect 139301 78099 139367 78102
rect 142110 78160 150131 78162
rect 142110 78104 150070 78160
rect 150126 78104 150131 78160
rect 142110 78102 150131 78104
rect 131798 77964 131804 78028
rect 131868 78026 131874 78028
rect 142110 78026 142170 78102
rect 150065 78099 150131 78102
rect 151118 78100 151124 78164
rect 151188 78162 151194 78164
rect 151445 78162 151511 78165
rect 151188 78160 151511 78162
rect 151188 78104 151450 78160
rect 151506 78104 151511 78160
rect 151188 78102 151511 78104
rect 151188 78100 151194 78102
rect 151445 78099 151511 78102
rect 152958 78100 152964 78164
rect 153028 78162 153034 78164
rect 153101 78162 153167 78165
rect 156321 78164 156387 78165
rect 176009 78164 176075 78165
rect 156270 78162 156276 78164
rect 153028 78160 153167 78162
rect 153028 78104 153106 78160
rect 153162 78104 153167 78160
rect 153028 78102 153167 78104
rect 156230 78102 156276 78162
rect 156340 78160 156387 78164
rect 175958 78162 175964 78164
rect 156382 78104 156387 78160
rect 153028 78100 153034 78102
rect 153101 78099 153167 78102
rect 156270 78100 156276 78102
rect 156340 78100 156387 78104
rect 175918 78102 175964 78162
rect 176028 78160 176075 78164
rect 176070 78104 176075 78160
rect 175958 78100 175964 78102
rect 176028 78100 176075 78104
rect 176150 78162 176210 78238
rect 176326 78236 176332 78300
rect 176396 78298 176402 78300
rect 176837 78298 176903 78301
rect 176396 78296 176903 78298
rect 176396 78240 176842 78296
rect 176898 78240 176903 78296
rect 176396 78238 176903 78240
rect 176396 78236 176402 78238
rect 176837 78235 176903 78238
rect 177849 78298 177915 78301
rect 203701 78298 203767 78301
rect 177849 78296 203767 78298
rect 177849 78240 177854 78296
rect 177910 78240 203706 78296
rect 203762 78240 203767 78296
rect 177849 78238 203767 78240
rect 177849 78235 177915 78238
rect 203701 78235 203767 78238
rect 198958 78162 198964 78164
rect 176150 78102 198964 78162
rect 198958 78100 198964 78102
rect 199028 78100 199034 78164
rect 156321 78099 156387 78100
rect 176009 78099 176075 78100
rect 131868 77966 142170 78026
rect 131868 77964 131874 77966
rect 147438 77964 147444 78028
rect 147508 78026 147514 78028
rect 160553 78026 160619 78029
rect 147508 78024 160619 78026
rect 147508 77968 160558 78024
rect 160614 77968 160619 78024
rect 147508 77966 160619 77968
rect 147508 77964 147514 77966
rect 160553 77963 160619 77966
rect 166390 77964 166396 78028
rect 166460 78026 166466 78028
rect 166717 78026 166783 78029
rect 166460 78024 166783 78026
rect 166460 77968 166722 78024
rect 166778 77968 166783 78024
rect 166460 77966 166783 77968
rect 166460 77964 166466 77966
rect 166717 77963 166783 77966
rect 171317 78026 171383 78029
rect 204161 78026 204227 78029
rect 269757 78026 269823 78029
rect 171317 78024 186330 78026
rect 171317 77968 171322 78024
rect 171378 77968 186330 78024
rect 171317 77966 186330 77968
rect 171317 77963 171383 77966
rect 60733 77890 60799 77893
rect 135805 77890 135871 77893
rect 136030 77890 136036 77892
rect 60733 77888 122850 77890
rect 60733 77832 60738 77888
rect 60794 77832 122850 77888
rect 60733 77830 122850 77832
rect 60733 77827 60799 77830
rect 122790 77754 122850 77830
rect 135805 77888 136036 77890
rect 135805 77832 135810 77888
rect 135866 77832 136036 77888
rect 135805 77830 136036 77832
rect 135805 77827 135871 77830
rect 136030 77828 136036 77830
rect 136100 77828 136106 77892
rect 138197 77890 138263 77893
rect 149421 77890 149487 77893
rect 138197 77888 149487 77890
rect 138197 77832 138202 77888
rect 138258 77832 149426 77888
rect 149482 77832 149487 77888
rect 138197 77830 149487 77832
rect 138197 77827 138263 77830
rect 149421 77827 149487 77830
rect 152774 77828 152780 77892
rect 152844 77890 152850 77892
rect 152917 77890 152983 77893
rect 152844 77888 152983 77890
rect 152844 77832 152922 77888
rect 152978 77832 152983 77888
rect 152844 77830 152983 77832
rect 152844 77828 152850 77830
rect 152917 77827 152983 77830
rect 153694 77828 153700 77892
rect 153764 77890 153770 77892
rect 154113 77890 154179 77893
rect 153764 77888 154179 77890
rect 153764 77832 154118 77888
rect 154174 77832 154179 77888
rect 153764 77830 154179 77832
rect 153764 77828 153770 77830
rect 154113 77827 154179 77830
rect 155401 77890 155467 77893
rect 155534 77890 155540 77892
rect 155401 77888 155540 77890
rect 155401 77832 155406 77888
rect 155462 77832 155540 77888
rect 155401 77830 155540 77832
rect 155401 77827 155467 77830
rect 155534 77828 155540 77830
rect 155604 77828 155610 77892
rect 156505 77890 156571 77893
rect 157006 77890 157012 77892
rect 156505 77888 157012 77890
rect 156505 77832 156510 77888
rect 156566 77832 157012 77888
rect 156505 77830 157012 77832
rect 156505 77827 156571 77830
rect 157006 77828 157012 77830
rect 157076 77828 157082 77892
rect 158294 77828 158300 77892
rect 158364 77890 158370 77892
rect 158621 77890 158687 77893
rect 158364 77888 158687 77890
rect 158364 77832 158626 77888
rect 158682 77832 158687 77888
rect 158364 77830 158687 77832
rect 158364 77828 158370 77830
rect 158621 77827 158687 77830
rect 171961 77890 172027 77893
rect 177062 77890 177068 77892
rect 171961 77888 177068 77890
rect 171961 77832 171966 77888
rect 172022 77832 177068 77888
rect 171961 77830 177068 77832
rect 171961 77827 172027 77830
rect 177062 77828 177068 77830
rect 177132 77828 177138 77892
rect 177205 77890 177271 77893
rect 179229 77890 179295 77893
rect 181529 77890 181595 77893
rect 177205 77888 181595 77890
rect 177205 77832 177210 77888
rect 177266 77832 179234 77888
rect 179290 77832 181534 77888
rect 181590 77832 181595 77888
rect 177205 77830 181595 77832
rect 177205 77827 177271 77830
rect 179229 77827 179295 77830
rect 181529 77827 181595 77830
rect 136909 77754 136975 77757
rect 122790 77752 136975 77754
rect 122790 77696 136914 77752
rect 136970 77696 136975 77752
rect 122790 77694 136975 77696
rect 136909 77691 136975 77694
rect 138013 77754 138079 77757
rect 138606 77754 138612 77756
rect 138013 77752 138612 77754
rect 138013 77696 138018 77752
rect 138074 77696 138612 77752
rect 138013 77694 138612 77696
rect 138013 77691 138079 77694
rect 138606 77692 138612 77694
rect 138676 77692 138682 77756
rect 139761 77754 139827 77757
rect 140630 77754 140636 77756
rect 139761 77752 140636 77754
rect 139761 77696 139766 77752
rect 139822 77696 140636 77752
rect 139761 77694 140636 77696
rect 139761 77691 139827 77694
rect 140630 77692 140636 77694
rect 140700 77692 140706 77756
rect 148409 77754 148475 77757
rect 148542 77754 148548 77756
rect 148409 77752 148548 77754
rect 148409 77696 148414 77752
rect 148470 77696 148548 77752
rect 148409 77694 148548 77696
rect 148409 77691 148475 77694
rect 148542 77692 148548 77694
rect 148612 77692 148618 77756
rect 149462 77692 149468 77756
rect 149532 77754 149538 77756
rect 157425 77754 157491 77757
rect 149532 77752 157491 77754
rect 149532 77696 157430 77752
rect 157486 77696 157491 77752
rect 149532 77694 157491 77696
rect 149532 77692 149538 77694
rect 157425 77691 157491 77694
rect 168557 77754 168623 77757
rect 168557 77752 173910 77754
rect 168557 77696 168562 77752
rect 168618 77696 173910 77752
rect 168557 77694 173910 77696
rect 168557 77691 168623 77694
rect 126462 77556 126468 77620
rect 126532 77618 126538 77620
rect 126532 77558 138030 77618
rect 126532 77556 126538 77558
rect 130326 77420 130332 77484
rect 130396 77482 130402 77484
rect 134057 77482 134123 77485
rect 130396 77480 134123 77482
rect 130396 77424 134062 77480
rect 134118 77424 134123 77480
rect 130396 77422 134123 77424
rect 137970 77482 138030 77558
rect 138238 77556 138244 77620
rect 138308 77618 138314 77620
rect 138749 77618 138815 77621
rect 138308 77616 138815 77618
rect 138308 77560 138754 77616
rect 138810 77560 138815 77616
rect 138308 77558 138815 77560
rect 138308 77556 138314 77558
rect 138749 77555 138815 77558
rect 139301 77618 139367 77621
rect 146937 77618 147003 77621
rect 153101 77618 153167 77621
rect 139301 77616 153167 77618
rect 139301 77560 139306 77616
rect 139362 77560 146942 77616
rect 146998 77560 153106 77616
rect 153162 77560 153167 77616
rect 139301 77558 153167 77560
rect 139301 77555 139367 77558
rect 146937 77555 147003 77558
rect 153101 77555 153167 77558
rect 156321 77618 156387 77621
rect 165061 77620 165127 77621
rect 156454 77618 156460 77620
rect 156321 77616 156460 77618
rect 156321 77560 156326 77616
rect 156382 77560 156460 77616
rect 156321 77558 156460 77560
rect 156321 77555 156387 77558
rect 156454 77556 156460 77558
rect 156524 77556 156530 77620
rect 165061 77616 165108 77620
rect 165172 77618 165178 77620
rect 170765 77618 170831 77621
rect 170990 77618 170996 77620
rect 165061 77560 165066 77616
rect 165061 77556 165108 77560
rect 165172 77558 165218 77618
rect 170765 77616 170996 77618
rect 170765 77560 170770 77616
rect 170826 77560 170996 77616
rect 170765 77558 170996 77560
rect 165172 77556 165178 77558
rect 165061 77555 165127 77556
rect 170765 77555 170831 77558
rect 170990 77556 170996 77558
rect 171060 77556 171066 77620
rect 171726 77556 171732 77620
rect 171796 77618 171802 77620
rect 172053 77618 172119 77621
rect 171796 77616 172119 77618
rect 171796 77560 172058 77616
rect 172114 77560 172119 77616
rect 171796 77558 172119 77560
rect 171796 77556 171802 77558
rect 172053 77555 172119 77558
rect 138105 77482 138171 77485
rect 137970 77480 138171 77482
rect 137970 77424 138110 77480
rect 138166 77424 138171 77480
rect 137970 77422 138171 77424
rect 130396 77420 130402 77422
rect 134057 77419 134123 77422
rect 138105 77419 138171 77422
rect 138289 77482 138355 77485
rect 140865 77484 140931 77485
rect 139158 77482 139164 77484
rect 138289 77480 139164 77482
rect 138289 77424 138294 77480
rect 138350 77424 139164 77480
rect 138289 77422 139164 77424
rect 138289 77419 138355 77422
rect 139158 77420 139164 77422
rect 139228 77420 139234 77484
rect 140814 77482 140820 77484
rect 140774 77422 140820 77482
rect 140884 77482 140931 77484
rect 141969 77482 142035 77485
rect 140884 77480 142035 77482
rect 140926 77424 141974 77480
rect 142030 77424 142035 77480
rect 140814 77420 140820 77422
rect 140884 77422 142035 77424
rect 173850 77482 173910 77694
rect 174486 77556 174492 77620
rect 174556 77618 174562 77620
rect 178033 77618 178099 77621
rect 174556 77616 178099 77618
rect 174556 77560 178038 77616
rect 178094 77560 178099 77616
rect 174556 77558 178099 77560
rect 174556 77556 174562 77558
rect 178033 77555 178099 77558
rect 182081 77482 182147 77485
rect 185577 77482 185643 77485
rect 173850 77422 176210 77482
rect 140884 77420 140931 77422
rect 140865 77419 140931 77420
rect 141969 77419 142035 77422
rect 134742 77346 134748 77348
rect 125550 77286 134748 77346
rect 100753 77210 100819 77213
rect 101581 77210 101647 77213
rect 125550 77210 125610 77286
rect 134742 77284 134748 77286
rect 134812 77284 134818 77348
rect 137553 77346 137619 77349
rect 138197 77346 138263 77349
rect 137553 77344 138263 77346
rect 137553 77288 137558 77344
rect 137614 77288 138202 77344
rect 138258 77288 138263 77344
rect 137553 77286 138263 77288
rect 137553 77283 137619 77286
rect 138197 77283 138263 77286
rect 139577 77346 139643 77349
rect 160829 77348 160895 77349
rect 161105 77348 161171 77349
rect 140262 77346 140268 77348
rect 139577 77344 140268 77346
rect 139577 77288 139582 77344
rect 139638 77288 140268 77344
rect 139577 77286 140268 77288
rect 139577 77283 139643 77286
rect 140262 77284 140268 77286
rect 140332 77284 140338 77348
rect 140814 77284 140820 77348
rect 140884 77346 140890 77348
rect 160829 77346 160876 77348
rect 140884 77286 141250 77346
rect 160784 77344 160876 77346
rect 160784 77288 160834 77344
rect 160784 77286 160876 77288
rect 140884 77284 140890 77286
rect 100753 77208 125610 77210
rect 100753 77152 100758 77208
rect 100814 77152 101586 77208
rect 101642 77152 125610 77208
rect 100753 77150 125610 77152
rect 134517 77210 134583 77213
rect 134926 77210 134932 77212
rect 134517 77208 134932 77210
rect 134517 77152 134522 77208
rect 134578 77152 134932 77208
rect 134517 77150 134932 77152
rect 100753 77147 100819 77150
rect 101581 77147 101647 77150
rect 134517 77147 134583 77150
rect 134926 77148 134932 77150
rect 134996 77148 135002 77212
rect 141190 77210 141250 77286
rect 160829 77284 160876 77286
rect 160940 77284 160946 77348
rect 161054 77284 161060 77348
rect 161124 77346 161171 77348
rect 176150 77346 176210 77422
rect 182081 77480 185643 77482
rect 182081 77424 182086 77480
rect 182142 77424 185582 77480
rect 185638 77424 185643 77480
rect 182081 77422 185643 77424
rect 186270 77482 186330 77966
rect 204161 78024 269823 78026
rect 204161 77968 204166 78024
rect 204222 77968 269762 78024
rect 269818 77968 269823 78024
rect 204161 77966 269823 77968
rect 204161 77963 204227 77966
rect 269757 77963 269823 77966
rect 187918 77828 187924 77892
rect 187988 77890 187994 77892
rect 287697 77890 287763 77893
rect 187988 77888 287763 77890
rect 187988 77832 287702 77888
rect 287758 77832 287763 77888
rect 187988 77830 287763 77832
rect 187988 77828 187994 77830
rect 287697 77827 287763 77830
rect 187693 77482 187759 77485
rect 186270 77480 187759 77482
rect 186270 77424 187698 77480
rect 187754 77424 187759 77480
rect 186270 77422 187759 77424
rect 182081 77419 182147 77422
rect 185577 77419 185643 77422
rect 187693 77419 187759 77422
rect 203149 77346 203215 77349
rect 204161 77346 204227 77349
rect 161124 77344 161216 77346
rect 161166 77288 161216 77344
rect 161124 77286 161216 77288
rect 176150 77344 204227 77346
rect 176150 77288 203154 77344
rect 203210 77288 204166 77344
rect 204222 77288 204227 77344
rect 176150 77286 204227 77288
rect 161124 77284 161171 77286
rect 160829 77283 160895 77284
rect 161105 77283 161171 77284
rect 203149 77283 203215 77286
rect 204161 77283 204227 77286
rect 141325 77210 141391 77213
rect 141190 77208 141391 77210
rect 141190 77152 141330 77208
rect 141386 77152 141391 77208
rect 141190 77150 141391 77152
rect 141325 77147 141391 77150
rect 142613 77210 142679 77213
rect 143022 77210 143028 77212
rect 142613 77208 143028 77210
rect 142613 77152 142618 77208
rect 142674 77152 143028 77208
rect 142613 77150 143028 77152
rect 142613 77147 142679 77150
rect 143022 77148 143028 77150
rect 143092 77148 143098 77212
rect 176142 77148 176148 77212
rect 176212 77210 176218 77212
rect 176285 77210 176351 77213
rect 176212 77208 176351 77210
rect 176212 77152 176290 77208
rect 176346 77152 176351 77208
rect 176212 77150 176351 77152
rect 176212 77148 176218 77150
rect 176285 77147 176351 77150
rect 178902 77148 178908 77212
rect 178972 77210 178978 77212
rect 179321 77210 179387 77213
rect 180057 77212 180123 77213
rect 180006 77210 180012 77212
rect 178972 77208 179387 77210
rect 178972 77152 179326 77208
rect 179382 77152 179387 77208
rect 178972 77150 179387 77152
rect 179966 77150 180012 77210
rect 180076 77208 180123 77212
rect 180118 77152 180123 77208
rect 178972 77148 178978 77150
rect 179321 77147 179387 77150
rect 180006 77148 180012 77150
rect 180076 77148 180123 77152
rect 180057 77147 180123 77148
rect 115657 77074 115723 77077
rect 146886 77074 146892 77076
rect 115657 77072 146892 77074
rect 115657 77016 115662 77072
rect 115718 77016 146892 77072
rect 115657 77014 146892 77016
rect 115657 77011 115723 77014
rect 146886 77012 146892 77014
rect 146956 77074 146962 77076
rect 147673 77074 147739 77077
rect 146956 77072 147739 77074
rect 146956 77016 147678 77072
rect 147734 77016 147739 77072
rect 146956 77014 147739 77016
rect 146956 77012 146962 77014
rect 147673 77011 147739 77014
rect 175089 77074 175155 77077
rect 191966 77074 191972 77076
rect 175089 77072 191972 77074
rect 175089 77016 175094 77072
rect 175150 77016 191972 77072
rect 175089 77014 191972 77016
rect 175089 77011 175155 77014
rect 191966 77012 191972 77014
rect 192036 77012 192042 77076
rect 117037 76938 117103 76941
rect 147305 76938 147371 76941
rect 154573 76938 154639 76941
rect 117037 76936 154639 76938
rect 117037 76880 117042 76936
rect 117098 76880 147310 76936
rect 147366 76880 154578 76936
rect 154634 76880 154639 76936
rect 117037 76878 154639 76880
rect 117037 76875 117103 76878
rect 147305 76875 147371 76878
rect 154573 76875 154639 76878
rect 169109 76938 169175 76941
rect 169334 76938 169340 76940
rect 169109 76936 169340 76938
rect 169109 76880 169114 76936
rect 169170 76880 169340 76936
rect 169109 76878 169340 76880
rect 169109 76875 169175 76878
rect 169334 76876 169340 76878
rect 169404 76876 169410 76940
rect 174854 76876 174860 76940
rect 174924 76938 174930 76940
rect 174997 76938 175063 76941
rect 174924 76936 175063 76938
rect 174924 76880 175002 76936
rect 175058 76880 175063 76936
rect 174924 76878 175063 76880
rect 174924 76876 174930 76878
rect 174997 76875 175063 76878
rect 178585 76938 178651 76941
rect 205909 76938 205975 76941
rect 178585 76936 205975 76938
rect 178585 76880 178590 76936
rect 178646 76880 205914 76936
rect 205970 76880 205975 76936
rect 178585 76878 205975 76880
rect 178585 76875 178651 76878
rect 205909 76875 205975 76878
rect 121085 76802 121151 76805
rect 148174 76802 148180 76804
rect 121085 76800 148180 76802
rect 121085 76744 121090 76800
rect 121146 76744 148180 76800
rect 121085 76742 148180 76744
rect 121085 76739 121151 76742
rect 148174 76740 148180 76742
rect 148244 76740 148250 76804
rect 157057 76802 157123 76805
rect 178534 76802 178540 76804
rect 157057 76800 178540 76802
rect 157057 76744 157062 76800
rect 157118 76744 178540 76800
rect 157057 76742 178540 76744
rect 157057 76739 157123 76742
rect 178534 76740 178540 76742
rect 178604 76740 178610 76804
rect 211797 76802 211863 76805
rect 200070 76800 211863 76802
rect 200070 76744 211802 76800
rect 211858 76744 211863 76800
rect 200070 76742 211863 76744
rect 113725 76666 113791 76669
rect 133505 76666 133571 76669
rect 113725 76664 133571 76666
rect 113725 76608 113730 76664
rect 113786 76608 133510 76664
rect 133566 76608 133571 76664
rect 113725 76606 133571 76608
rect 113725 76603 113791 76606
rect 133505 76603 133571 76606
rect 134241 76666 134307 76669
rect 153929 76668 153995 76669
rect 134374 76666 134380 76668
rect 134241 76664 134380 76666
rect 134241 76608 134246 76664
rect 134302 76608 134380 76664
rect 134241 76606 134380 76608
rect 134241 76603 134307 76606
rect 134374 76604 134380 76606
rect 134444 76604 134450 76668
rect 153878 76666 153884 76668
rect 153838 76606 153884 76666
rect 153948 76664 153995 76668
rect 153990 76608 153995 76664
rect 153878 76604 153884 76606
rect 153948 76604 153995 76608
rect 170254 76604 170260 76668
rect 170324 76666 170330 76668
rect 170765 76666 170831 76669
rect 191598 76666 191604 76668
rect 170324 76664 191604 76666
rect 170324 76608 170770 76664
rect 170826 76608 191604 76664
rect 170324 76606 191604 76608
rect 170324 76604 170330 76606
rect 153929 76603 153995 76604
rect 170765 76603 170831 76606
rect 191598 76604 191604 76606
rect 191668 76604 191674 76668
rect 34513 76530 34579 76533
rect 100753 76530 100819 76533
rect 34513 76528 100819 76530
rect 34513 76472 34518 76528
rect 34574 76472 100758 76528
rect 100814 76472 100819 76528
rect 34513 76470 100819 76472
rect 34513 76467 34579 76470
rect 100753 76467 100819 76470
rect 130377 76530 130443 76533
rect 133597 76530 133663 76533
rect 130377 76528 133663 76530
rect 130377 76472 130382 76528
rect 130438 76472 133602 76528
rect 133658 76472 133663 76528
rect 130377 76470 133663 76472
rect 130377 76467 130443 76470
rect 133597 76467 133663 76470
rect 162301 76530 162367 76533
rect 162526 76530 162532 76532
rect 162301 76528 162532 76530
rect 162301 76472 162306 76528
rect 162362 76472 162532 76528
rect 162301 76470 162532 76472
rect 162301 76467 162367 76470
rect 162526 76468 162532 76470
rect 162596 76468 162602 76532
rect 170213 76530 170279 76533
rect 170806 76530 170812 76532
rect 170213 76528 170812 76530
rect 170213 76472 170218 76528
rect 170274 76472 170812 76528
rect 170213 76470 170812 76472
rect 170213 76467 170279 76470
rect 170806 76468 170812 76470
rect 170876 76468 170882 76532
rect 171593 76530 171659 76533
rect 186681 76530 186747 76533
rect 171593 76528 186747 76530
rect 171593 76472 171598 76528
rect 171654 76472 186686 76528
rect 186742 76472 186747 76528
rect 171593 76470 186747 76472
rect 171593 76467 171659 76470
rect 186681 76467 186747 76470
rect 130285 76394 130351 76397
rect 134057 76394 134123 76397
rect 130285 76392 134123 76394
rect 130285 76336 130290 76392
rect 130346 76336 134062 76392
rect 134118 76336 134123 76392
rect 130285 76334 134123 76336
rect 130285 76331 130351 76334
rect 134057 76331 134123 76334
rect 151629 76394 151695 76397
rect 183686 76394 183692 76396
rect 151629 76392 183692 76394
rect 151629 76336 151634 76392
rect 151690 76336 183692 76392
rect 151629 76334 183692 76336
rect 151629 76331 151695 76334
rect 183686 76332 183692 76334
rect 183756 76394 183762 76396
rect 200070 76394 200130 76742
rect 211797 76739 211863 76742
rect 204621 76666 204687 76669
rect 247677 76666 247743 76669
rect 204621 76664 247743 76666
rect 204621 76608 204626 76664
rect 204682 76608 247682 76664
rect 247738 76608 247743 76664
rect 204621 76606 247743 76608
rect 204621 76603 204687 76606
rect 183756 76334 200130 76394
rect 183756 76332 183762 76334
rect 152825 76258 152891 76261
rect 204854 76258 204914 76606
rect 247677 76603 247743 76606
rect 205909 76530 205975 76533
rect 553393 76530 553459 76533
rect 205909 76528 553459 76530
rect 205909 76472 205914 76528
rect 205970 76472 553398 76528
rect 553454 76472 553459 76528
rect 205909 76470 553459 76472
rect 205909 76467 205975 76470
rect 553393 76467 553459 76470
rect 152825 76256 204914 76258
rect 152825 76200 152830 76256
rect 152886 76200 204914 76256
rect 152825 76198 204914 76200
rect 152825 76195 152891 76198
rect 163313 76124 163379 76125
rect 163262 76122 163268 76124
rect 163222 76062 163268 76122
rect 163332 76120 163379 76124
rect 163374 76064 163379 76120
rect 163262 76060 163268 76062
rect 163332 76060 163379 76064
rect 163313 76059 163379 76060
rect 164969 76122 165035 76125
rect 165470 76122 165476 76124
rect 164969 76120 165476 76122
rect 164969 76064 164974 76120
rect 165030 76064 165476 76120
rect 164969 76062 165476 76064
rect 164969 76059 165035 76062
rect 165470 76060 165476 76062
rect 165540 76060 165546 76124
rect 130377 75986 130443 75989
rect 131665 75986 131731 75989
rect 130377 75984 131731 75986
rect 130377 75928 130382 75984
rect 130438 75928 131670 75984
rect 131726 75928 131731 75984
rect 130377 75926 131731 75928
rect 130377 75923 130443 75926
rect 131665 75923 131731 75926
rect 134006 75924 134012 75988
rect 134076 75986 134082 75988
rect 134701 75986 134767 75989
rect 134076 75984 134767 75986
rect 134076 75928 134706 75984
rect 134762 75928 134767 75984
rect 134076 75926 134767 75928
rect 134076 75924 134082 75926
rect 134701 75923 134767 75926
rect 135437 75986 135503 75989
rect 135897 75988 135963 75989
rect 135662 75986 135668 75988
rect 135437 75984 135668 75986
rect 135437 75928 135442 75984
rect 135498 75928 135668 75984
rect 135437 75926 135668 75928
rect 135437 75923 135503 75926
rect 135662 75924 135668 75926
rect 135732 75924 135738 75988
rect 135846 75924 135852 75988
rect 135916 75986 135963 75988
rect 148133 75986 148199 75989
rect 148726 75986 148732 75988
rect 135916 75984 136008 75986
rect 135958 75928 136008 75984
rect 135916 75926 136008 75928
rect 148133 75984 148732 75986
rect 148133 75928 148138 75984
rect 148194 75928 148732 75984
rect 148133 75926 148732 75928
rect 135916 75924 135963 75926
rect 135897 75923 135963 75924
rect 148133 75923 148199 75926
rect 148726 75924 148732 75926
rect 148796 75924 148802 75988
rect 162577 75986 162643 75989
rect 162710 75986 162716 75988
rect 162577 75984 162716 75986
rect 162577 75928 162582 75984
rect 162638 75928 162716 75984
rect 162577 75926 162716 75928
rect 162577 75923 162643 75926
rect 162710 75924 162716 75926
rect 162780 75924 162786 75988
rect 163446 75924 163452 75988
rect 163516 75986 163522 75988
rect 163681 75986 163747 75989
rect 166441 75988 166507 75989
rect 166390 75986 166396 75988
rect 163516 75984 163747 75986
rect 163516 75928 163686 75984
rect 163742 75928 163747 75984
rect 163516 75926 163747 75928
rect 166350 75926 166396 75986
rect 166460 75984 166507 75988
rect 166502 75928 166507 75984
rect 163516 75924 163522 75926
rect 163681 75923 163747 75926
rect 166390 75924 166396 75926
rect 166460 75924 166507 75928
rect 166574 75924 166580 75988
rect 166644 75986 166650 75988
rect 166809 75986 166875 75989
rect 166644 75984 166875 75986
rect 166644 75928 166814 75984
rect 166870 75928 166875 75984
rect 166644 75926 166875 75928
rect 166644 75924 166650 75926
rect 166441 75923 166507 75924
rect 166809 75923 166875 75926
rect 167678 75924 167684 75988
rect 167748 75986 167754 75988
rect 168189 75986 168255 75989
rect 167748 75984 168255 75986
rect 167748 75928 168194 75984
rect 168250 75928 168255 75984
rect 167748 75926 168255 75928
rect 167748 75924 167754 75926
rect 168189 75923 168255 75926
rect 173566 75924 173572 75988
rect 173636 75986 173642 75988
rect 173801 75986 173867 75989
rect 173636 75984 173867 75986
rect 173636 75928 173806 75984
rect 173862 75928 173867 75984
rect 173636 75926 173867 75928
rect 173636 75924 173642 75926
rect 173801 75923 173867 75926
rect 119521 75850 119587 75853
rect 129733 75850 129799 75853
rect 131021 75850 131087 75853
rect 119521 75848 131087 75850
rect 119521 75792 119526 75848
rect 119582 75792 129738 75848
rect 129794 75792 131026 75848
rect 131082 75792 131087 75848
rect 119521 75790 131087 75792
rect 119521 75787 119587 75790
rect 129733 75787 129799 75790
rect 131021 75787 131087 75790
rect 135345 75850 135411 75853
rect 135478 75850 135484 75852
rect 135345 75848 135484 75850
rect 135345 75792 135350 75848
rect 135406 75792 135484 75848
rect 135345 75790 135484 75792
rect 135345 75787 135411 75790
rect 135478 75788 135484 75790
rect 135548 75788 135554 75852
rect 187325 75850 187391 75853
rect 157290 75848 187391 75850
rect 157290 75792 187330 75848
rect 187386 75792 187391 75848
rect 157290 75790 187391 75792
rect 106733 75714 106799 75717
rect 139342 75714 139348 75716
rect 103470 75712 139348 75714
rect 103470 75656 106738 75712
rect 106794 75656 139348 75712
rect 103470 75654 139348 75656
rect 96613 75170 96679 75173
rect 103470 75170 103530 75654
rect 106733 75651 106799 75654
rect 139342 75652 139348 75654
rect 139412 75652 139418 75716
rect 152958 75652 152964 75716
rect 153028 75714 153034 75716
rect 157290 75714 157350 75790
rect 187325 75787 187391 75790
rect 153028 75654 157350 75714
rect 174077 75714 174143 75717
rect 206185 75714 206251 75717
rect 206553 75714 206619 75717
rect 174077 75712 206619 75714
rect 174077 75656 174082 75712
rect 174138 75656 206190 75712
rect 206246 75656 206558 75712
rect 206614 75656 206619 75712
rect 174077 75654 206619 75656
rect 153028 75652 153034 75654
rect 174077 75651 174143 75654
rect 206185 75651 206251 75654
rect 206553 75651 206619 75654
rect 110965 75578 111031 75581
rect 174721 75580 174787 75581
rect 140998 75578 141004 75580
rect 110965 75576 141004 75578
rect 110965 75520 110970 75576
rect 111026 75520 141004 75576
rect 110965 75518 141004 75520
rect 110965 75515 111031 75518
rect 140998 75516 141004 75518
rect 141068 75516 141074 75580
rect 174670 75578 174676 75580
rect 174630 75518 174676 75578
rect 174740 75576 174787 75580
rect 174782 75520 174787 75576
rect 174670 75516 174676 75518
rect 174740 75516 174787 75520
rect 175590 75516 175596 75580
rect 175660 75578 175666 75580
rect 176561 75578 176627 75581
rect 193254 75578 193260 75580
rect 175660 75576 193260 75578
rect 175660 75520 176566 75576
rect 176622 75520 193260 75576
rect 175660 75518 193260 75520
rect 175660 75516 175666 75518
rect 174721 75515 174787 75516
rect 176561 75515 176627 75518
rect 193254 75516 193260 75518
rect 193324 75516 193330 75580
rect 121177 75442 121243 75445
rect 145598 75442 145604 75444
rect 121177 75440 145604 75442
rect 121177 75384 121182 75440
rect 121238 75384 145604 75440
rect 121177 75382 145604 75384
rect 121177 75379 121243 75382
rect 145598 75380 145604 75382
rect 145668 75442 145674 75444
rect 145925 75442 145991 75445
rect 145668 75440 145991 75442
rect 145668 75384 145930 75440
rect 145986 75384 145991 75440
rect 145668 75382 145991 75384
rect 145668 75380 145674 75382
rect 145925 75379 145991 75382
rect 174537 75442 174603 75445
rect 174721 75442 174787 75445
rect 196382 75442 196388 75444
rect 174537 75440 196388 75442
rect 174537 75384 174542 75440
rect 174598 75384 174726 75440
rect 174782 75384 196388 75440
rect 174537 75382 196388 75384
rect 174537 75379 174603 75382
rect 174721 75379 174787 75382
rect 196382 75380 196388 75382
rect 196452 75380 196458 75444
rect 122649 75306 122715 75309
rect 146109 75306 146175 75309
rect 157425 75306 157491 75309
rect 122649 75304 157491 75306
rect 122649 75248 122654 75304
rect 122710 75248 146114 75304
rect 146170 75248 157430 75304
rect 157486 75248 157491 75304
rect 122649 75246 157491 75248
rect 122649 75243 122715 75246
rect 146109 75243 146175 75246
rect 157425 75243 157491 75246
rect 171174 75244 171180 75308
rect 171244 75306 171250 75308
rect 453297 75306 453363 75309
rect 171244 75304 453363 75306
rect 171244 75248 453302 75304
rect 453358 75248 453363 75304
rect 171244 75246 453363 75248
rect 171244 75244 171250 75246
rect 453297 75243 453363 75246
rect 96613 75168 103530 75170
rect 96613 75112 96618 75168
rect 96674 75112 103530 75168
rect 96613 75110 103530 75112
rect 121913 75170 121979 75173
rect 144729 75170 144795 75173
rect 121913 75168 144795 75170
rect 121913 75112 121918 75168
rect 121974 75112 144734 75168
rect 144790 75112 144795 75168
rect 121913 75110 144795 75112
rect 96613 75107 96679 75110
rect 121913 75107 121979 75110
rect 144729 75107 144795 75110
rect 170990 75108 170996 75172
rect 171060 75170 171066 75172
rect 188061 75170 188127 75173
rect 171060 75168 188127 75170
rect 171060 75112 188066 75168
rect 188122 75112 188127 75168
rect 171060 75110 188127 75112
rect 171060 75108 171066 75110
rect 188061 75107 188127 75110
rect 206553 75170 206619 75173
rect 535453 75170 535519 75173
rect 206553 75168 535519 75170
rect 206553 75112 206558 75168
rect 206614 75112 535458 75168
rect 535514 75112 535519 75168
rect 206553 75110 535519 75112
rect 206553 75107 206619 75110
rect 535453 75107 535519 75110
rect 115749 75034 115815 75037
rect 148358 75034 148364 75036
rect 115749 75032 148364 75034
rect 115749 74976 115754 75032
rect 115810 74976 148364 75032
rect 115749 74974 148364 74976
rect 115749 74971 115815 74974
rect 148358 74972 148364 74974
rect 148428 74972 148434 75036
rect 155309 75034 155375 75037
rect 181110 75034 181116 75036
rect 155309 75032 181116 75034
rect 155309 74976 155314 75032
rect 155370 74976 181116 75032
rect 155309 74974 181116 74976
rect 155309 74971 155375 74974
rect 181110 74972 181116 74974
rect 181180 74972 181186 75036
rect 183553 75034 183619 75037
rect 189022 75034 189028 75036
rect 183553 75032 189028 75034
rect 183553 74976 183558 75032
rect 183614 74976 189028 75032
rect 183553 74974 189028 74976
rect 183553 74971 183619 74974
rect 189022 74972 189028 74974
rect 189092 74972 189098 75036
rect 136725 74898 136791 74901
rect 137502 74898 137508 74900
rect 136725 74896 137508 74898
rect 136725 74840 136730 74896
rect 136786 74840 137508 74896
rect 136725 74838 137508 74840
rect 136725 74835 136791 74838
rect 137502 74836 137508 74838
rect 137572 74836 137578 74900
rect 144545 74762 144611 74765
rect 144678 74762 144684 74764
rect 144545 74760 144684 74762
rect 144545 74704 144550 74760
rect 144606 74704 144684 74760
rect 144545 74702 144684 74704
rect 144545 74699 144611 74702
rect 144678 74700 144684 74702
rect 144748 74700 144754 74764
rect 122465 74626 122531 74629
rect 122782 74626 122788 74628
rect 122465 74624 122788 74626
rect 122465 74568 122470 74624
rect 122526 74568 122788 74624
rect 122465 74566 122788 74568
rect 122465 74563 122531 74566
rect 122782 74564 122788 74566
rect 122852 74564 122858 74628
rect 118550 74428 118556 74492
rect 118620 74490 118626 74492
rect 152273 74490 152339 74493
rect 118620 74488 152339 74490
rect 118620 74432 152278 74488
rect 152334 74432 152339 74488
rect 118620 74430 152339 74432
rect 118620 74428 118626 74430
rect 152273 74427 152339 74430
rect 156454 74428 156460 74492
rect 156524 74490 156530 74492
rect 191465 74490 191531 74493
rect 156524 74488 191531 74490
rect 156524 74432 191470 74488
rect 191526 74432 191531 74488
rect 156524 74430 191531 74432
rect 156524 74428 156530 74430
rect 191465 74427 191531 74430
rect 122782 74292 122788 74356
rect 122852 74354 122858 74356
rect 157977 74354 158043 74357
rect 158253 74354 158319 74357
rect 122852 74352 158319 74354
rect 122852 74296 157982 74352
rect 158038 74296 158258 74352
rect 158314 74296 158319 74352
rect 122852 74294 158319 74296
rect 122852 74292 122858 74294
rect 157977 74291 158043 74294
rect 158253 74291 158319 74294
rect 173893 74354 173959 74357
rect 174905 74354 174971 74357
rect 193806 74354 193812 74356
rect 173893 74352 193812 74354
rect 173893 74296 173898 74352
rect 173954 74296 174910 74352
rect 174966 74296 193812 74352
rect 173893 74294 193812 74296
rect 173893 74291 173959 74294
rect 174905 74291 174971 74294
rect 193806 74292 193812 74294
rect 193876 74292 193882 74356
rect 134149 74218 134215 74221
rect 134374 74218 134380 74220
rect 134149 74216 134380 74218
rect 134149 74160 134154 74216
rect 134210 74160 134380 74216
rect 134149 74158 134380 74160
rect 134149 74155 134215 74158
rect 134374 74156 134380 74158
rect 134444 74156 134450 74220
rect 155677 74218 155743 74221
rect 183502 74218 183508 74220
rect 155677 74216 183508 74218
rect 155677 74160 155682 74216
rect 155738 74160 183508 74216
rect 155677 74158 183508 74160
rect 155677 74155 155743 74158
rect 183502 74156 183508 74158
rect 183572 74156 183578 74220
rect 112529 74082 112595 74085
rect 139710 74082 139716 74084
rect 112529 74080 139716 74082
rect 112529 74024 112534 74080
rect 112590 74024 139716 74080
rect 112529 74022 139716 74024
rect 112529 74019 112595 74022
rect 139710 74020 139716 74022
rect 139780 74020 139786 74084
rect 158069 74082 158135 74085
rect 158621 74082 158687 74085
rect 158069 74080 158687 74082
rect 158069 74024 158074 74080
rect 158130 74024 158626 74080
rect 158682 74024 158687 74080
rect 158069 74022 158687 74024
rect 158069 74019 158135 74022
rect 158621 74019 158687 74022
rect 177062 74020 177068 74084
rect 177132 74082 177138 74084
rect 187734 74082 187740 74084
rect 177132 74022 187740 74082
rect 177132 74020 177138 74022
rect 187734 74020 187740 74022
rect 187804 74020 187810 74084
rect 114921 73946 114987 73949
rect 140814 73946 140820 73948
rect 114921 73944 140820 73946
rect 114921 73888 114926 73944
rect 114982 73888 140820 73944
rect 114921 73886 140820 73888
rect 114921 73883 114987 73886
rect 140814 73884 140820 73886
rect 140884 73884 140890 73948
rect 145046 73884 145052 73948
rect 145116 73946 145122 73948
rect 145833 73946 145899 73949
rect 145116 73944 145899 73946
rect 145116 73888 145838 73944
rect 145894 73888 145899 73944
rect 145116 73886 145899 73888
rect 145116 73884 145122 73886
rect 145833 73883 145899 73886
rect 175181 73946 175247 73949
rect 175457 73946 175523 73949
rect 192518 73946 192524 73948
rect 175181 73944 192524 73946
rect 175181 73888 175186 73944
rect 175242 73888 175462 73944
rect 175518 73888 192524 73944
rect 175181 73886 192524 73888
rect 175181 73883 175247 73886
rect 175457 73883 175523 73886
rect 192518 73884 192524 73886
rect 192588 73884 192594 73948
rect 122598 73748 122604 73812
rect 122668 73810 122674 73812
rect 155309 73810 155375 73813
rect 122668 73808 155375 73810
rect 122668 73752 155314 73808
rect 155370 73752 155375 73808
rect 122668 73750 155375 73752
rect 122668 73748 122674 73750
rect 155309 73747 155375 73750
rect 158621 73810 158687 73813
rect 181294 73810 181300 73812
rect 158621 73808 181300 73810
rect 158621 73752 158626 73808
rect 158682 73752 181300 73808
rect 158621 73750 181300 73752
rect 158621 73747 158687 73750
rect 181294 73748 181300 73750
rect 181364 73748 181370 73812
rect 191465 73810 191531 73813
rect 304993 73810 305059 73813
rect 191465 73808 305059 73810
rect 191465 73752 191470 73808
rect 191526 73752 304998 73808
rect 305054 73752 305059 73808
rect 191465 73750 305059 73752
rect 191465 73747 191531 73750
rect 304993 73747 305059 73750
rect 152273 73674 152339 73677
rect 152733 73674 152799 73677
rect 152273 73672 152799 73674
rect 152273 73616 152278 73672
rect 152334 73616 152738 73672
rect 152794 73616 152799 73672
rect 152273 73614 152799 73616
rect 152273 73611 152339 73614
rect 152733 73611 152799 73614
rect 158478 73612 158484 73676
rect 158548 73674 158554 73676
rect 179822 73674 179828 73676
rect 158548 73614 179828 73674
rect 158548 73612 158554 73614
rect 179822 73612 179828 73614
rect 179892 73612 179898 73676
rect 122414 73068 122420 73132
rect 122484 73130 122490 73132
rect 156321 73130 156387 73133
rect 122484 73128 156387 73130
rect 122484 73072 156326 73128
rect 156382 73072 156387 73128
rect 122484 73070 156387 73072
rect 122484 73068 122490 73070
rect 156321 73067 156387 73070
rect 156822 73068 156828 73132
rect 156892 73130 156898 73132
rect 205633 73130 205699 73133
rect 156892 73128 205699 73130
rect 156892 73072 205638 73128
rect 205694 73072 205699 73128
rect 156892 73070 205699 73072
rect 156892 73068 156898 73070
rect 205633 73067 205699 73070
rect 105629 72994 105695 72997
rect 139526 72994 139532 72996
rect 105629 72992 139532 72994
rect 105629 72936 105634 72992
rect 105690 72936 139532 72992
rect 105629 72934 139532 72936
rect 105629 72931 105695 72934
rect 139526 72932 139532 72934
rect 139596 72932 139602 72996
rect 155953 72994 156019 72997
rect 157149 72994 157215 72997
rect 183134 72994 183140 72996
rect 155953 72992 183140 72994
rect 155953 72936 155958 72992
rect 156014 72936 157154 72992
rect 157210 72936 183140 72992
rect 155953 72934 183140 72936
rect 155953 72931 156019 72934
rect 157149 72931 157215 72934
rect 183134 72932 183140 72934
rect 183204 72932 183210 72996
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 118601 72858 118667 72861
rect 151118 72858 151124 72860
rect 118601 72856 151124 72858
rect 118601 72800 118606 72856
rect 118662 72800 151124 72856
rect 118601 72798 151124 72800
rect 118601 72795 118667 72798
rect 151118 72796 151124 72798
rect 151188 72796 151194 72860
rect 175641 72858 175707 72861
rect 176469 72858 176535 72861
rect 196566 72858 196572 72860
rect 175641 72856 196572 72858
rect 175641 72800 175646 72856
rect 175702 72800 176474 72856
rect 176530 72800 196572 72856
rect 175641 72798 196572 72800
rect 175641 72795 175707 72798
rect 176469 72795 176535 72798
rect 196566 72796 196572 72798
rect 196636 72796 196642 72860
rect 583520 72844 584960 72934
rect 117129 72722 117195 72725
rect 149094 72722 149100 72724
rect 117129 72720 149100 72722
rect 117129 72664 117134 72720
rect 117190 72664 149100 72720
rect 117129 72662 149100 72664
rect 117129 72659 117195 72662
rect 149094 72660 149100 72662
rect 149164 72722 149170 72724
rect 149462 72722 149468 72724
rect 149164 72662 149468 72722
rect 149164 72660 149170 72662
rect 149462 72660 149468 72662
rect 149532 72660 149538 72724
rect 123845 72586 123911 72589
rect 150014 72586 150020 72588
rect 123845 72584 150020 72586
rect 123845 72528 123850 72584
rect 123906 72528 150020 72584
rect 123845 72526 150020 72528
rect 123845 72523 123911 72526
rect 150014 72524 150020 72526
rect 150084 72524 150090 72588
rect 157425 72450 157491 72453
rect 178033 72450 178099 72453
rect 157425 72448 178099 72450
rect 157425 72392 157430 72448
rect 157486 72392 178038 72448
rect 178094 72392 178099 72448
rect 157425 72390 178099 72392
rect 157425 72387 157491 72390
rect 178033 72387 178099 72390
rect 205633 72450 205699 72453
rect 301497 72450 301563 72453
rect 205633 72448 301563 72450
rect 205633 72392 205638 72448
rect 205694 72392 301502 72448
rect 301558 72392 301563 72448
rect 205633 72390 301563 72392
rect 205633 72387 205699 72390
rect 301497 72387 301563 72390
rect 145414 72252 145420 72316
rect 145484 72314 145490 72316
rect 156597 72314 156663 72317
rect 145484 72312 156663 72314
rect 145484 72256 156602 72312
rect 156658 72256 156663 72312
rect 145484 72254 156663 72256
rect 145484 72252 145490 72254
rect 156597 72251 156663 72254
rect 116301 71770 116367 71773
rect 156873 71770 156939 71773
rect 116301 71768 156939 71770
rect -960 71634 480 71724
rect 116301 71712 116306 71768
rect 116362 71712 156878 71768
rect 156934 71712 156939 71768
rect 116301 71710 156939 71712
rect 116301 71707 116367 71710
rect 156873 71707 156939 71710
rect 159817 71770 159883 71773
rect 184974 71770 184980 71772
rect 159817 71768 184980 71770
rect 159817 71712 159822 71768
rect 159878 71712 184980 71768
rect 159817 71710 184980 71712
rect 159817 71707 159883 71710
rect 184974 71708 184980 71710
rect 185044 71708 185050 71772
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 118182 71572 118188 71636
rect 118252 71634 118258 71636
rect 152406 71634 152412 71636
rect 118252 71574 152412 71634
rect 118252 71572 118258 71574
rect 152406 71572 152412 71574
rect 152476 71572 152482 71636
rect 173566 71572 173572 71636
rect 173636 71634 173642 71636
rect 197486 71634 197492 71636
rect 173636 71574 197492 71634
rect 173636 71572 173642 71574
rect 197486 71572 197492 71574
rect 197556 71572 197562 71636
rect 116761 71498 116827 71501
rect 149646 71498 149652 71500
rect 116761 71496 149652 71498
rect 116761 71440 116766 71496
rect 116822 71440 149652 71496
rect 116761 71438 149652 71440
rect 116761 71435 116827 71438
rect 149646 71436 149652 71438
rect 149716 71436 149722 71500
rect 164049 71498 164115 71501
rect 184054 71498 184060 71500
rect 164049 71496 184060 71498
rect 164049 71440 164054 71496
rect 164110 71440 184060 71496
rect 164049 71438 184060 71440
rect 164049 71435 164115 71438
rect 184054 71436 184060 71438
rect 184124 71436 184130 71500
rect 114461 71362 114527 71365
rect 145046 71362 145052 71364
rect 114461 71360 145052 71362
rect 114461 71304 114466 71360
rect 114522 71304 145052 71360
rect 114461 71302 145052 71304
rect 114461 71299 114527 71302
rect 145046 71300 145052 71302
rect 145116 71300 145122 71364
rect 188429 71362 188495 71365
rect 489177 71362 489243 71365
rect 188429 71360 489243 71362
rect 188429 71304 188434 71360
rect 188490 71304 489182 71360
rect 489238 71304 489243 71360
rect 188429 71302 489243 71304
rect 188429 71299 188495 71302
rect 489177 71299 489243 71302
rect 187734 71164 187740 71228
rect 187804 71226 187810 71228
rect 507853 71226 507919 71229
rect 187804 71224 507919 71226
rect 187804 71168 507858 71224
rect 507914 71168 507919 71224
rect 187804 71166 507919 71168
rect 187804 71164 187810 71166
rect 507853 71163 507919 71166
rect 144126 71028 144132 71092
rect 144196 71090 144202 71092
rect 144729 71090 144795 71093
rect 144196 71088 144795 71090
rect 144196 71032 144734 71088
rect 144790 71032 144795 71088
rect 144196 71030 144795 71032
rect 144196 71028 144202 71030
rect 144729 71027 144795 71030
rect 197486 71028 197492 71092
rect 197556 71090 197562 71092
rect 198038 71090 198044 71092
rect 197556 71030 198044 71090
rect 197556 71028 197562 71030
rect 198038 71028 198044 71030
rect 198108 71090 198114 71092
rect 531313 71090 531379 71093
rect 198108 71088 531379 71090
rect 198108 71032 531318 71088
rect 531374 71032 531379 71088
rect 198108 71030 531379 71032
rect 198108 71028 198114 71030
rect 531313 71027 531379 71030
rect 142061 70412 142127 70413
rect 142061 70408 142108 70412
rect 142172 70410 142178 70412
rect 142061 70352 142066 70408
rect 142061 70348 142108 70352
rect 142172 70350 142218 70410
rect 142172 70348 142178 70350
rect 142061 70347 142127 70348
rect 122230 70212 122236 70276
rect 122300 70274 122306 70276
rect 156045 70274 156111 70277
rect 122300 70272 156111 70274
rect 122300 70216 156050 70272
rect 156106 70216 156111 70272
rect 122300 70214 156111 70216
rect 122300 70212 122306 70214
rect 156045 70211 156111 70214
rect 175958 70212 175964 70276
rect 176028 70274 176034 70276
rect 201350 70274 201356 70276
rect 176028 70214 201356 70274
rect 176028 70212 176034 70214
rect 201350 70212 201356 70214
rect 201420 70212 201426 70276
rect 128905 70138 128971 70141
rect 103470 70136 128971 70138
rect 103470 70080 128910 70136
rect 128966 70080 128971 70136
rect 103470 70078 128971 70080
rect 41413 69594 41479 69597
rect 102869 69594 102935 69597
rect 103470 69594 103530 70078
rect 128905 70075 128971 70078
rect 148726 70076 148732 70140
rect 148796 70138 148802 70140
rect 182766 70138 182772 70140
rect 148796 70078 182772 70138
rect 148796 70076 148802 70078
rect 182766 70076 182772 70078
rect 182836 70138 182842 70140
rect 182836 70078 184674 70138
rect 182836 70076 182842 70078
rect 115105 70002 115171 70005
rect 144494 70002 144500 70004
rect 115105 70000 144500 70002
rect 115105 69944 115110 70000
rect 115166 69944 144500 70000
rect 115105 69942 144500 69944
rect 115105 69939 115171 69942
rect 144494 69940 144500 69942
rect 144564 69940 144570 70004
rect 147213 70002 147279 70005
rect 178350 70002 178356 70004
rect 147213 70000 178356 70002
rect 147213 69944 147218 70000
rect 147274 69944 178356 70000
rect 147213 69942 178356 69944
rect 147213 69939 147279 69942
rect 178350 69940 178356 69942
rect 178420 70002 178426 70004
rect 182909 70002 182975 70005
rect 178420 70000 182975 70002
rect 178420 69944 182914 70000
rect 182970 69944 182975 70000
rect 178420 69942 182975 69944
rect 178420 69940 178426 69942
rect 182909 69939 182975 69942
rect 156045 69866 156111 69869
rect 156781 69866 156847 69869
rect 156045 69864 156847 69866
rect 156045 69808 156050 69864
rect 156106 69808 156786 69864
rect 156842 69808 156847 69864
rect 156045 69806 156847 69808
rect 156045 69803 156111 69806
rect 156781 69803 156847 69806
rect 41413 69592 103530 69594
rect 41413 69536 41418 69592
rect 41474 69536 102874 69592
rect 102930 69536 103530 69592
rect 41413 69534 103530 69536
rect 184614 69594 184674 70078
rect 187417 69730 187483 69733
rect 498193 69730 498259 69733
rect 187417 69728 498259 69730
rect 187417 69672 187422 69728
rect 187478 69672 498198 69728
rect 498254 69672 498259 69728
rect 187417 69670 498259 69672
rect 187417 69667 187483 69670
rect 498193 69667 498259 69670
rect 200757 69594 200823 69597
rect 184614 69592 200823 69594
rect 184614 69536 200762 69592
rect 200818 69536 200823 69592
rect 184614 69534 200823 69536
rect 41413 69531 41479 69534
rect 102869 69531 102935 69534
rect 200757 69531 200823 69534
rect 201350 69532 201356 69596
rect 201420 69594 201426 69596
rect 561673 69594 561739 69597
rect 201420 69592 561739 69594
rect 201420 69536 561678 69592
rect 561734 69536 561739 69592
rect 201420 69534 561739 69536
rect 201420 69532 201426 69534
rect 561673 69531 561739 69534
rect 114369 68914 114435 68917
rect 144678 68914 144684 68916
rect 114369 68912 144684 68914
rect 114369 68856 114374 68912
rect 114430 68856 144684 68912
rect 114369 68854 144684 68856
rect 114369 68851 114435 68854
rect 144678 68852 144684 68854
rect 144748 68852 144754 68916
rect 145598 68852 145604 68916
rect 145668 68914 145674 68916
rect 148317 68914 148383 68917
rect 183001 68916 183067 68917
rect 182950 68914 182956 68916
rect 145668 68912 148383 68914
rect 145668 68856 148322 68912
rect 148378 68856 148383 68912
rect 145668 68854 148383 68856
rect 182910 68854 182956 68914
rect 183020 68912 183067 68916
rect 183062 68856 183067 68912
rect 145668 68852 145674 68854
rect 148317 68851 148383 68854
rect 182950 68852 182956 68854
rect 183020 68852 183067 68856
rect 198774 68852 198780 68916
rect 198844 68914 198850 68916
rect 199377 68914 199443 68917
rect 198844 68912 199443 68914
rect 198844 68856 199382 68912
rect 199438 68856 199443 68912
rect 198844 68854 199443 68856
rect 198844 68852 198850 68854
rect 183001 68851 183067 68852
rect 199377 68851 199443 68854
rect 114829 68778 114895 68781
rect 114829 68776 122850 68778
rect 114829 68720 114834 68776
rect 114890 68720 122850 68776
rect 114829 68718 122850 68720
rect 114829 68715 114895 68718
rect 122790 68642 122850 68718
rect 176142 68716 176148 68780
rect 176212 68778 176218 68780
rect 176212 68718 200130 68778
rect 176212 68716 176218 68718
rect 144310 68642 144316 68644
rect 122790 68582 144316 68642
rect 144310 68580 144316 68582
rect 144380 68580 144386 68644
rect 148542 68308 148548 68372
rect 148612 68370 148618 68372
rect 184197 68370 184263 68373
rect 148612 68368 184263 68370
rect 148612 68312 184202 68368
rect 184258 68312 184263 68368
rect 148612 68310 184263 68312
rect 148612 68308 148618 68310
rect 184197 68307 184263 68310
rect 8937 68234 9003 68237
rect 132217 68234 132283 68237
rect 8937 68232 132283 68234
rect 8937 68176 8942 68232
rect 8998 68176 132222 68232
rect 132278 68176 132283 68232
rect 8937 68174 132283 68176
rect 8937 68171 9003 68174
rect 132217 68171 132283 68174
rect 154573 68234 154639 68237
rect 189717 68234 189783 68237
rect 154573 68232 189783 68234
rect 154573 68176 154578 68232
rect 154634 68176 189722 68232
rect 189778 68176 189783 68232
rect 154573 68174 189783 68176
rect 200070 68234 200130 68718
rect 203609 68234 203675 68237
rect 565813 68234 565879 68237
rect 200070 68232 565879 68234
rect 200070 68176 203614 68232
rect 203670 68176 565818 68232
rect 565874 68176 565879 68232
rect 200070 68174 565879 68176
rect 154573 68171 154639 68174
rect 189717 68171 189783 68174
rect 203609 68171 203675 68174
rect 565813 68171 565879 68174
rect 104249 67554 104315 67557
rect 135662 67554 135668 67556
rect 103470 67552 135668 67554
rect 103470 67496 104254 67552
rect 104310 67496 135668 67552
rect 103470 67494 135668 67496
rect 40033 67010 40099 67013
rect 103470 67010 103530 67494
rect 104249 67491 104315 67494
rect 135662 67492 135668 67494
rect 135732 67492 135738 67556
rect 189022 67492 189028 67556
rect 189092 67554 189098 67556
rect 189165 67554 189231 67557
rect 189092 67552 189231 67554
rect 189092 67496 189170 67552
rect 189226 67496 189231 67552
rect 189092 67494 189231 67496
rect 189092 67492 189098 67494
rect 189165 67491 189231 67494
rect 155534 67356 155540 67420
rect 155604 67418 155610 67420
rect 189349 67418 189415 67421
rect 189901 67418 189967 67421
rect 155604 67416 189967 67418
rect 155604 67360 189354 67416
rect 189410 67360 189906 67416
rect 189962 67360 189967 67416
rect 155604 67358 189967 67360
rect 155604 67356 155610 67358
rect 189349 67355 189415 67358
rect 189901 67355 189967 67358
rect 151486 67220 151492 67284
rect 151556 67282 151562 67284
rect 178166 67282 178172 67284
rect 151556 67222 178172 67282
rect 151556 67220 151562 67222
rect 178166 67220 178172 67222
rect 178236 67282 178242 67284
rect 242893 67282 242959 67285
rect 178236 67280 242959 67282
rect 178236 67224 242898 67280
rect 242954 67224 242959 67280
rect 178236 67222 242959 67224
rect 178236 67220 178242 67222
rect 242893 67219 242959 67222
rect 148174 67084 148180 67148
rect 148244 67146 148250 67148
rect 213913 67146 213979 67149
rect 148244 67144 213979 67146
rect 148244 67088 213918 67144
rect 213974 67088 213979 67144
rect 148244 67086 213979 67088
rect 148244 67084 148250 67086
rect 213913 67083 213979 67086
rect 40033 67008 103530 67010
rect 40033 66952 40038 67008
rect 40094 66952 103530 67008
rect 40033 66950 103530 66952
rect 189901 67010 189967 67013
rect 295333 67010 295399 67013
rect 189901 67008 295399 67010
rect 189901 66952 189906 67008
rect 189962 66952 295338 67008
rect 295394 66952 295399 67008
rect 189901 66950 295399 66952
rect 40033 66947 40099 66950
rect 189901 66947 189967 66950
rect 295333 66947 295399 66950
rect 11053 66874 11119 66877
rect 133638 66874 133644 66876
rect 11053 66872 133644 66874
rect 11053 66816 11058 66872
rect 11114 66816 133644 66872
rect 11053 66814 133644 66816
rect 11053 66811 11119 66814
rect 133638 66812 133644 66814
rect 133708 66812 133714 66876
rect 146886 66812 146892 66876
rect 146956 66874 146962 66876
rect 193857 66874 193923 66877
rect 376753 66874 376819 66877
rect 146956 66872 193923 66874
rect 146956 66816 193862 66872
rect 193918 66816 193923 66872
rect 146956 66814 193923 66816
rect 146956 66812 146962 66814
rect 193857 66811 193923 66814
rect 200070 66872 376819 66874
rect 200070 66816 376758 66872
rect 376814 66816 376819 66872
rect 200070 66814 376819 66816
rect 162158 66676 162164 66740
rect 162228 66738 162234 66740
rect 196157 66738 196223 66741
rect 200070 66738 200130 66814
rect 376753 66811 376819 66814
rect 162228 66736 200130 66738
rect 162228 66680 196162 66736
rect 196218 66680 200130 66736
rect 162228 66678 200130 66680
rect 162228 66676 162234 66678
rect 196157 66675 196223 66678
rect 105445 66194 105511 66197
rect 106181 66194 106247 66197
rect 137502 66194 137508 66196
rect 105445 66192 137508 66194
rect 105445 66136 105450 66192
rect 105506 66136 106186 66192
rect 106242 66136 137508 66192
rect 105445 66134 137508 66136
rect 105445 66131 105511 66134
rect 106181 66131 106247 66134
rect 137502 66132 137508 66134
rect 137572 66132 137578 66196
rect 153878 66132 153884 66196
rect 153948 66194 153954 66196
rect 187877 66194 187943 66197
rect 153948 66192 187943 66194
rect 153948 66136 187882 66192
rect 187938 66136 187943 66192
rect 153948 66134 187943 66136
rect 153948 66132 153954 66134
rect 187877 66131 187943 66134
rect 160686 65996 160692 66060
rect 160756 66058 160762 66060
rect 193581 66058 193647 66061
rect 194501 66058 194567 66061
rect 160756 66056 194567 66058
rect 160756 66000 193586 66056
rect 193642 66000 194506 66056
rect 194562 66000 194567 66056
rect 160756 65998 194567 66000
rect 160756 65996 160762 65998
rect 193581 65995 193647 65998
rect 194501 65995 194567 65998
rect 187877 65922 187943 65925
rect 274633 65922 274699 65925
rect 187877 65920 274699 65922
rect 187877 65864 187882 65920
rect 187938 65864 274638 65920
rect 274694 65864 274699 65920
rect 187877 65862 274699 65864
rect 187877 65859 187943 65862
rect 274633 65859 274699 65862
rect 171910 65724 171916 65788
rect 171980 65786 171986 65788
rect 189390 65786 189396 65788
rect 171980 65726 189396 65786
rect 171980 65724 171986 65726
rect 189390 65724 189396 65726
rect 189460 65786 189466 65788
rect 194501 65786 194567 65789
rect 362953 65786 363019 65789
rect 189460 65726 190470 65786
rect 189460 65724 189466 65726
rect 190410 65650 190470 65726
rect 194501 65784 363019 65786
rect 194501 65728 194506 65784
rect 194562 65728 362958 65784
rect 363014 65728 363019 65784
rect 194501 65726 363019 65728
rect 194501 65723 194567 65726
rect 362953 65723 363019 65726
rect 514017 65650 514083 65653
rect 190410 65648 514083 65650
rect 190410 65592 514022 65648
rect 514078 65592 514083 65648
rect 190410 65590 514083 65592
rect 514017 65587 514083 65590
rect 57237 65514 57303 65517
rect 105445 65514 105511 65517
rect 57237 65512 105511 65514
rect 57237 65456 57242 65512
rect 57298 65456 105450 65512
rect 105506 65456 105511 65512
rect 57237 65454 105511 65456
rect 57237 65451 57303 65454
rect 105445 65451 105511 65454
rect 173750 65452 173756 65516
rect 173820 65514 173826 65516
rect 195094 65514 195100 65516
rect 173820 65454 195100 65514
rect 173820 65452 173826 65454
rect 195094 65452 195100 65454
rect 195164 65514 195170 65516
rect 527817 65514 527883 65517
rect 195164 65512 527883 65514
rect 195164 65456 527822 65512
rect 527878 65456 527883 65512
rect 195164 65454 527883 65456
rect 195164 65452 195170 65454
rect 527817 65451 527883 65454
rect 142061 64972 142127 64973
rect 142061 64970 142108 64972
rect 142016 64968 142108 64970
rect 142172 64970 142178 64972
rect 142016 64912 142066 64968
rect 142016 64910 142108 64912
rect 142061 64908 142108 64910
rect 142172 64910 142254 64970
rect 142172 64908 142178 64910
rect 142061 64907 142127 64908
rect 142061 64834 142127 64837
rect 142016 64832 142170 64834
rect 142016 64776 142066 64832
rect 142122 64776 142170 64832
rect 142016 64774 142170 64776
rect 142061 64771 142170 64774
rect 174670 64772 174676 64836
rect 174740 64834 174746 64836
rect 197854 64834 197860 64836
rect 174740 64774 197860 64834
rect 174740 64772 174746 64774
rect 197854 64772 197860 64774
rect 197924 64772 197930 64836
rect 142110 64700 142170 64771
rect 142102 64636 142108 64700
rect 142172 64636 142178 64700
rect 172094 64636 172100 64700
rect 172164 64698 172170 64700
rect 186998 64698 187004 64700
rect 172164 64638 187004 64698
rect 172164 64636 172170 64638
rect 186998 64636 187004 64638
rect 187068 64636 187074 64700
rect 186998 64228 187004 64292
rect 187068 64290 187074 64292
rect 511993 64290 512059 64293
rect 187068 64288 512059 64290
rect 187068 64232 511998 64288
rect 512054 64232 512059 64288
rect 187068 64230 512059 64232
rect 187068 64228 187074 64230
rect 511993 64227 512059 64230
rect 197854 64092 197860 64156
rect 197924 64154 197930 64156
rect 543733 64154 543799 64157
rect 197924 64152 543799 64154
rect 197924 64096 543738 64152
rect 543794 64096 543799 64152
rect 197924 64094 543799 64096
rect 197924 64092 197930 64094
rect 543733 64091 543799 64094
rect 110413 63474 110479 63477
rect 111701 63474 111767 63477
rect 138606 63474 138612 63476
rect 110413 63472 138612 63474
rect 110413 63416 110418 63472
rect 110474 63416 111706 63472
rect 111762 63416 138612 63472
rect 110413 63414 138612 63416
rect 110413 63411 110479 63414
rect 111701 63411 111767 63414
rect 138606 63412 138612 63414
rect 138676 63412 138682 63476
rect 166206 63412 166212 63476
rect 166276 63474 166282 63476
rect 200297 63474 200363 63477
rect 201401 63474 201467 63477
rect 166276 63472 201467 63474
rect 166276 63416 200302 63472
rect 200358 63416 201406 63472
rect 201462 63416 201467 63472
rect 166276 63414 201467 63416
rect 166276 63412 166282 63414
rect 200297 63411 200363 63414
rect 201401 63411 201467 63414
rect 149462 63276 149468 63340
rect 149532 63338 149538 63340
rect 227713 63338 227779 63341
rect 149532 63336 227779 63338
rect 149532 63280 227718 63336
rect 227774 63280 227779 63336
rect 149532 63278 227779 63280
rect 149532 63276 149538 63278
rect 227713 63275 227779 63278
rect 154062 63140 154068 63204
rect 154132 63202 154138 63204
rect 187785 63202 187851 63205
rect 277393 63202 277459 63205
rect 154132 63200 277459 63202
rect 154132 63144 187790 63200
rect 187846 63144 277398 63200
rect 277454 63144 277459 63200
rect 154132 63142 277459 63144
rect 154132 63140 154138 63142
rect 187785 63139 187851 63142
rect 277393 63139 277459 63142
rect 155718 63004 155724 63068
rect 155788 63066 155794 63068
rect 189073 63066 189139 63069
rect 292573 63066 292639 63069
rect 155788 63064 292639 63066
rect 155788 63008 189078 63064
rect 189134 63008 292578 63064
rect 292634 63008 292639 63064
rect 155788 63006 292639 63008
rect 155788 63004 155794 63006
rect 189073 63003 189139 63006
rect 292573 63003 292639 63006
rect 174854 62868 174860 62932
rect 174924 62930 174930 62932
rect 197302 62930 197308 62932
rect 174924 62870 197308 62930
rect 174924 62868 174930 62870
rect 197302 62868 197308 62870
rect 197372 62930 197378 62932
rect 201401 62930 201467 62933
rect 430573 62930 430639 62933
rect 197372 62870 200130 62930
rect 197372 62868 197378 62870
rect 75177 62794 75243 62797
rect 110413 62794 110479 62797
rect 75177 62792 110479 62794
rect 75177 62736 75182 62792
rect 75238 62736 110418 62792
rect 110474 62736 110479 62792
rect 75177 62734 110479 62736
rect 200070 62794 200130 62870
rect 201401 62928 430639 62930
rect 201401 62872 201406 62928
rect 201462 62872 430578 62928
rect 430634 62872 430639 62928
rect 201401 62870 430639 62872
rect 201401 62867 201467 62870
rect 430573 62867 430639 62870
rect 547873 62794 547939 62797
rect 200070 62792 547939 62794
rect 200070 62736 547878 62792
rect 547934 62736 547939 62792
rect 200070 62734 547939 62736
rect 75177 62731 75243 62734
rect 110413 62731 110479 62734
rect 547873 62731 547939 62734
rect 186957 62114 187023 62117
rect 196065 62116 196131 62117
rect 187182 62114 187188 62116
rect 186957 62112 187188 62114
rect 186957 62056 186962 62112
rect 187018 62056 187188 62112
rect 186957 62054 187188 62056
rect 186957 62051 187023 62054
rect 187182 62052 187188 62054
rect 187252 62052 187258 62116
rect 196014 62114 196020 62116
rect 195974 62054 196020 62114
rect 196084 62112 196131 62116
rect 196126 62056 196131 62112
rect 196014 62052 196020 62054
rect 196084 62052 196131 62056
rect 196065 62051 196131 62052
rect 157006 61916 157012 61980
rect 157076 61978 157082 61980
rect 190637 61978 190703 61981
rect 191741 61978 191807 61981
rect 157076 61976 191807 61978
rect 157076 61920 190642 61976
rect 190698 61920 191746 61976
rect 191802 61920 191807 61976
rect 157076 61918 191807 61920
rect 157076 61916 157082 61918
rect 190637 61915 190703 61918
rect 191741 61915 191807 61918
rect 164918 61780 164924 61844
rect 164988 61842 164994 61844
rect 199009 61842 199075 61845
rect 164988 61840 199075 61842
rect 164988 61784 199014 61840
rect 199070 61784 199075 61840
rect 164988 61782 199075 61784
rect 164988 61780 164994 61782
rect 199009 61779 199075 61782
rect 149830 61644 149836 61708
rect 149900 61706 149906 61708
rect 231853 61706 231919 61709
rect 149900 61704 231919 61706
rect 149900 61648 231858 61704
rect 231914 61648 231919 61704
rect 149900 61646 231919 61648
rect 149900 61644 149906 61646
rect 231853 61643 231919 61646
rect 191741 61570 191807 61573
rect 309133 61570 309199 61573
rect 191741 61568 309199 61570
rect 191741 61512 191746 61568
rect 191802 61512 309138 61568
rect 309194 61512 309199 61568
rect 191741 61510 309199 61512
rect 191741 61507 191807 61510
rect 309133 61507 309199 61510
rect 199009 61434 199075 61437
rect 422937 61434 423003 61437
rect 199009 61432 423003 61434
rect 199009 61376 199014 61432
rect 199070 61376 422942 61432
rect 422998 61376 423003 61432
rect 199009 61374 423003 61376
rect 199009 61371 199075 61374
rect 422937 61371 423003 61374
rect 165102 60556 165108 60620
rect 165172 60618 165178 60620
rect 198917 60618 198983 60621
rect 165172 60616 200130 60618
rect 165172 60560 198922 60616
rect 198978 60560 200130 60616
rect 165172 60558 200130 60560
rect 165172 60556 165178 60558
rect 198917 60555 198983 60558
rect 176326 60420 176332 60484
rect 176396 60482 176402 60484
rect 176396 60422 180810 60482
rect 176396 60420 176402 60422
rect 180750 59938 180810 60422
rect 200070 60074 200130 60558
rect 412633 60074 412699 60077
rect 200070 60072 412699 60074
rect 200070 60016 412638 60072
rect 412694 60016 412699 60072
rect 200070 60014 412699 60016
rect 412633 60011 412699 60014
rect 200982 59938 200988 59940
rect 180750 59878 200988 59938
rect 200982 59876 200988 59878
rect 201052 59938 201058 59940
rect 567837 59938 567903 59941
rect 201052 59936 567903 59938
rect 201052 59880 567842 59936
rect 567898 59880 567903 59936
rect 201052 59878 567903 59880
rect 201052 59876 201058 59878
rect 567837 59875 567903 59878
rect 583520 59666 584960 59756
rect 567150 59606 584960 59666
rect 188286 59332 188292 59396
rect 188356 59394 188362 59396
rect 567150 59394 567210 59606
rect 583520 59516 584960 59606
rect 188356 59334 567210 59394
rect 188356 59332 188362 59334
rect 167494 59196 167500 59260
rect 167564 59258 167570 59260
rect 201861 59258 201927 59261
rect 202781 59258 202847 59261
rect 167564 59256 202847 59258
rect 167564 59200 201866 59256
rect 201922 59200 202786 59256
rect 202842 59200 202847 59256
rect 167564 59198 202847 59200
rect 167564 59196 167570 59198
rect 201861 59195 201927 59198
rect 202781 59195 202847 59198
rect 154246 59060 154252 59124
rect 154316 59122 154322 59124
rect 188245 59122 188311 59125
rect 154316 59120 190470 59122
rect 154316 59064 188250 59120
rect 188306 59064 190470 59120
rect 154316 59062 190470 59064
rect 154316 59060 154322 59062
rect 188245 59059 188311 59062
rect 190410 58986 190470 59062
rect 281533 58986 281599 58989
rect 190410 58984 281599 58986
rect 190410 58928 281538 58984
rect 281594 58928 281599 58984
rect 190410 58926 281599 58928
rect 281533 58923 281599 58926
rect 157926 58788 157932 58852
rect 157996 58850 158002 58852
rect 191925 58850 191991 58853
rect 327073 58850 327139 58853
rect 157996 58848 327139 58850
rect 157996 58792 191930 58848
rect 191986 58792 327078 58848
rect 327134 58792 327139 58848
rect 157996 58790 327139 58792
rect 157996 58788 158002 58790
rect 191925 58787 191991 58790
rect 327073 58787 327139 58790
rect -960 58578 480 58668
rect 162342 58652 162348 58716
rect 162412 58714 162418 58716
rect 196157 58714 196223 58717
rect 380893 58714 380959 58717
rect 162412 58712 380959 58714
rect 162412 58656 196162 58712
rect 196218 58656 380898 58712
rect 380954 58656 380959 58712
rect 162412 58654 380959 58656
rect 162412 58652 162418 58654
rect 196157 58651 196223 58654
rect 380893 58651 380959 58654
rect 202781 58578 202847 58581
rect 450537 58578 450603 58581
rect -960 58518 674 58578
rect -960 58442 480 58518
rect 614 58442 674 58518
rect 202781 58576 450603 58578
rect 202781 58520 202786 58576
rect 202842 58520 450542 58576
rect 450598 58520 450603 58576
rect 202781 58518 450603 58520
rect 202781 58515 202847 58518
rect 450537 58515 450603 58518
rect -960 58428 674 58442
rect 246 58382 674 58428
rect 246 58034 306 58382
rect 120758 58034 120764 58036
rect 246 57974 120764 58034
rect 120758 57972 120764 57974
rect 120828 57972 120834 58036
rect 100753 57898 100819 57901
rect 101673 57898 101739 57901
rect 134374 57898 134380 57900
rect 100753 57896 134380 57898
rect 100753 57840 100758 57896
rect 100814 57840 101678 57896
rect 101734 57840 134380 57896
rect 100753 57838 134380 57840
rect 100753 57835 100819 57838
rect 101673 57835 101739 57838
rect 134374 57836 134380 57838
rect 134444 57836 134450 57900
rect 152774 57836 152780 57900
rect 152844 57898 152850 57900
rect 186589 57898 186655 57901
rect 152844 57896 190470 57898
rect 152844 57840 186594 57896
rect 186650 57840 190470 57896
rect 152844 57838 190470 57840
rect 152844 57836 152850 57838
rect 186589 57835 186655 57838
rect 138422 57762 138428 57764
rect 113130 57702 138428 57762
rect 77293 57354 77359 57357
rect 110321 57354 110387 57357
rect 113130 57354 113190 57702
rect 138422 57700 138428 57702
rect 138492 57700 138498 57764
rect 190410 57762 190470 57838
rect 263593 57762 263659 57765
rect 190410 57760 263659 57762
rect 190410 57704 263598 57760
rect 263654 57704 263659 57760
rect 190410 57702 263659 57704
rect 263593 57699 263659 57702
rect 156638 57564 156644 57628
rect 156708 57626 156714 57628
rect 190545 57626 190611 57629
rect 313273 57626 313339 57629
rect 156708 57624 313339 57626
rect 156708 57568 190550 57624
rect 190606 57568 313278 57624
rect 313334 57568 313339 57624
rect 156708 57566 313339 57568
rect 156708 57564 156714 57566
rect 190545 57563 190611 57566
rect 313273 57563 313339 57566
rect 160870 57428 160876 57492
rect 160940 57490 160946 57492
rect 193765 57490 193831 57493
rect 364977 57490 365043 57493
rect 160940 57488 365043 57490
rect 160940 57432 193770 57488
rect 193826 57432 364982 57488
rect 365038 57432 365043 57488
rect 160940 57430 365043 57432
rect 160940 57428 160946 57430
rect 193765 57427 193831 57430
rect 364977 57427 365043 57430
rect 77293 57352 113190 57354
rect 77293 57296 77298 57352
rect 77354 57296 110326 57352
rect 110382 57296 113190 57352
rect 77293 57294 113190 57296
rect 77293 57291 77359 57294
rect 110321 57291 110387 57294
rect 165286 57292 165292 57356
rect 165356 57354 165362 57356
rect 198825 57354 198891 57357
rect 414657 57354 414723 57357
rect 165356 57352 414723 57354
rect 165356 57296 198830 57352
rect 198886 57296 414662 57352
rect 414718 57296 414723 57352
rect 165356 57294 414723 57296
rect 165356 57292 165362 57294
rect 198825 57291 198891 57294
rect 414657 57291 414723 57294
rect 25497 57218 25563 57221
rect 100753 57218 100819 57221
rect 25497 57216 100819 57218
rect 25497 57160 25502 57216
rect 25558 57160 100758 57216
rect 100814 57160 100819 57216
rect 25497 57158 100819 57160
rect 25497 57155 25563 57158
rect 100753 57155 100819 57158
rect 175038 57156 175044 57220
rect 175108 57218 175114 57220
rect 200798 57218 200804 57220
rect 175108 57158 200804 57218
rect 175108 57156 175114 57158
rect 200798 57156 200804 57158
rect 200868 57218 200874 57220
rect 545757 57218 545823 57221
rect 200868 57216 545823 57218
rect 200868 57160 545762 57216
rect 545818 57160 545823 57216
rect 200868 57158 545823 57160
rect 200868 57156 200874 57158
rect 545757 57155 545823 57158
rect 167678 56476 167684 56540
rect 167748 56538 167754 56540
rect 201953 56538 202019 56541
rect 202781 56538 202847 56541
rect 167748 56536 202847 56538
rect 167748 56480 201958 56536
rect 202014 56480 202786 56536
rect 202842 56480 202847 56536
rect 167748 56478 202847 56480
rect 167748 56476 167754 56478
rect 201953 56475 202019 56478
rect 202781 56475 202847 56478
rect 158846 56340 158852 56404
rect 158916 56402 158922 56404
rect 190821 56402 190887 56405
rect 349153 56402 349219 56405
rect 158916 56400 349219 56402
rect 158916 56344 190826 56400
rect 190882 56344 349158 56400
rect 349214 56344 349219 56400
rect 158916 56342 349219 56344
rect 158916 56340 158922 56342
rect 190821 56339 190887 56342
rect 349153 56339 349219 56342
rect 163262 56204 163268 56268
rect 163332 56266 163338 56268
rect 197353 56266 197419 56269
rect 398833 56266 398899 56269
rect 163332 56264 398899 56266
rect 163332 56208 197358 56264
rect 197414 56208 398838 56264
rect 398894 56208 398899 56264
rect 163332 56206 398899 56208
rect 163332 56204 163338 56206
rect 197353 56203 197419 56206
rect 398833 56203 398899 56206
rect 176510 56068 176516 56132
rect 176580 56130 176586 56132
rect 200614 56130 200620 56132
rect 176580 56070 200620 56130
rect 176580 56068 176586 56070
rect 200614 56068 200620 56070
rect 200684 56130 200690 56132
rect 201350 56130 201356 56132
rect 200684 56070 201356 56130
rect 200684 56068 200690 56070
rect 201350 56068 201356 56070
rect 201420 56068 201426 56132
rect 202781 56130 202847 56133
rect 459553 56130 459619 56133
rect 202781 56128 459619 56130
rect 202781 56072 202786 56128
rect 202842 56072 459558 56128
rect 459614 56072 459619 56128
rect 202781 56070 459619 56072
rect 202781 56067 202847 56070
rect 459553 56067 459619 56070
rect 172278 55932 172284 55996
rect 172348 55994 172354 55996
rect 204253 55994 204319 55997
rect 499573 55994 499639 55997
rect 172348 55992 499639 55994
rect 172348 55936 204258 55992
rect 204314 55936 499578 55992
rect 499634 55936 499639 55992
rect 172348 55934 499639 55936
rect 172348 55932 172354 55934
rect 204253 55931 204319 55934
rect 499573 55931 499639 55934
rect 201350 55796 201356 55860
rect 201420 55858 201426 55860
rect 563697 55858 563763 55861
rect 201420 55856 563763 55858
rect 201420 55800 563702 55856
rect 563758 55800 563763 55856
rect 201420 55798 563763 55800
rect 201420 55796 201426 55798
rect 563697 55795 563763 55798
rect 142061 55316 142127 55317
rect 142061 55314 142108 55316
rect 142016 55312 142108 55314
rect 142172 55314 142178 55316
rect 142016 55256 142066 55312
rect 142016 55254 142108 55256
rect 142061 55252 142108 55254
rect 142172 55254 142254 55314
rect 142172 55252 142178 55254
rect 142061 55251 142127 55252
rect 111793 55178 111859 55181
rect 113081 55178 113147 55181
rect 138238 55178 138244 55180
rect 111793 55176 138244 55178
rect 111793 55120 111798 55176
rect 111854 55120 113086 55176
rect 113142 55120 138244 55176
rect 111793 55118 138244 55120
rect 111793 55115 111859 55118
rect 113081 55115 113147 55118
rect 138238 55116 138244 55118
rect 138308 55116 138314 55180
rect 142061 55178 142127 55181
rect 142016 55176 142170 55178
rect 142016 55120 142066 55176
rect 142122 55120 142170 55176
rect 142016 55118 142170 55120
rect 142061 55115 142170 55118
rect 163446 55116 163452 55180
rect 163516 55178 163522 55180
rect 197445 55178 197511 55181
rect 163516 55176 197511 55178
rect 163516 55120 197450 55176
rect 197506 55120 197511 55176
rect 163516 55118 197511 55120
rect 163516 55116 163522 55118
rect 197445 55115 197511 55118
rect 201677 55180 201743 55181
rect 201677 55176 201724 55180
rect 201788 55178 201794 55180
rect 201677 55120 201682 55176
rect 201677 55116 201724 55120
rect 201788 55118 201834 55178
rect 201788 55116 201794 55118
rect 201677 55115 201743 55116
rect 142110 55044 142170 55115
rect 142102 54980 142108 55044
rect 142172 54980 142178 55044
rect 158110 54980 158116 55044
rect 158180 55042 158186 55044
rect 191833 55042 191899 55045
rect 158180 55040 191899 55042
rect 158180 54984 191838 55040
rect 191894 54984 191899 55040
rect 158180 54982 191899 54984
rect 158180 54980 158186 54982
rect 191833 54979 191899 54982
rect 161054 54844 161060 54908
rect 161124 54906 161130 54908
rect 193397 54906 193463 54909
rect 161124 54904 193463 54906
rect 161124 54848 193402 54904
rect 193458 54848 193463 54904
rect 161124 54846 193463 54848
rect 161124 54844 161130 54846
rect 193397 54843 193463 54846
rect 191833 54770 191899 54773
rect 331213 54770 331279 54773
rect 191833 54768 331279 54770
rect 191833 54712 191838 54768
rect 191894 54712 331218 54768
rect 331274 54712 331279 54768
rect 191833 54710 331279 54712
rect 191833 54707 191899 54710
rect 331213 54707 331279 54710
rect 193397 54634 193463 54637
rect 369853 54634 369919 54637
rect 193397 54632 369919 54634
rect 193397 54576 193402 54632
rect 193458 54576 369858 54632
rect 369914 54576 369919 54632
rect 193397 54574 369919 54576
rect 193397 54571 193463 54574
rect 369853 54571 369919 54574
rect 84193 54498 84259 54501
rect 111793 54498 111859 54501
rect 84193 54496 111859 54498
rect 84193 54440 84198 54496
rect 84254 54440 111798 54496
rect 111854 54440 111859 54496
rect 84193 54438 111859 54440
rect 84193 54435 84259 54438
rect 111793 54435 111859 54438
rect 197445 54498 197511 54501
rect 401593 54498 401659 54501
rect 197445 54496 401659 54498
rect 197445 54440 197450 54496
rect 197506 54440 401598 54496
rect 401654 54440 401659 54496
rect 197445 54438 401659 54440
rect 197445 54435 197511 54438
rect 401593 54435 401659 54438
rect 166390 53756 166396 53820
rect 166460 53818 166466 53820
rect 200205 53818 200271 53821
rect 201401 53818 201467 53821
rect 166460 53816 201467 53818
rect 166460 53760 200210 53816
rect 200266 53760 201406 53816
rect 201462 53760 201467 53816
rect 166460 53758 201467 53760
rect 166460 53756 166466 53758
rect 200205 53755 200271 53758
rect 201401 53755 201467 53758
rect 162526 53620 162532 53684
rect 162596 53682 162602 53684
rect 194777 53682 194843 53685
rect 162596 53680 194843 53682
rect 162596 53624 194782 53680
rect 194838 53624 194843 53680
rect 162596 53622 194843 53624
rect 162596 53620 162602 53622
rect 194777 53619 194843 53622
rect 154430 53484 154436 53548
rect 154500 53546 154506 53548
rect 154500 53486 180810 53546
rect 154500 53484 154506 53486
rect 180750 53410 180810 53486
rect 182582 53410 182588 53412
rect 180750 53350 182588 53410
rect 182582 53348 182588 53350
rect 182652 53410 182658 53412
rect 284385 53410 284451 53413
rect 182652 53408 284451 53410
rect 182652 53352 284390 53408
rect 284446 53352 284451 53408
rect 182652 53350 284451 53352
rect 182652 53348 182658 53350
rect 284385 53347 284451 53350
rect 194777 53274 194843 53277
rect 382917 53274 382983 53277
rect 194777 53272 382983 53274
rect 194777 53216 194782 53272
rect 194838 53216 382922 53272
rect 382978 53216 382983 53272
rect 194777 53214 382983 53216
rect 194777 53211 194843 53214
rect 382917 53211 382983 53214
rect 201401 53138 201467 53141
rect 437473 53138 437539 53141
rect 201401 53136 437539 53138
rect 201401 53080 201406 53136
rect 201462 53080 437478 53136
rect 437534 53080 437539 53136
rect 201401 53078 437539 53080
rect 201401 53075 201467 53078
rect 437473 53075 437539 53078
rect 100753 52458 100819 52461
rect 102041 52458 102107 52461
rect 134190 52458 134196 52460
rect 100753 52456 134196 52458
rect 100753 52400 100758 52456
rect 100814 52400 102046 52456
rect 102102 52400 134196 52456
rect 100753 52398 134196 52400
rect 100753 52395 100819 52398
rect 102041 52395 102107 52398
rect 134190 52396 134196 52398
rect 134260 52396 134266 52460
rect 167862 52396 167868 52460
rect 167932 52458 167938 52460
rect 201769 52458 201835 52461
rect 202781 52458 202847 52461
rect 167932 52456 202847 52458
rect 167932 52400 201774 52456
rect 201830 52400 202786 52456
rect 202842 52400 202847 52456
rect 167932 52398 202847 52400
rect 167932 52396 167938 52398
rect 201769 52395 201835 52398
rect 202781 52395 202847 52398
rect 163630 52260 163636 52324
rect 163700 52322 163706 52324
rect 194685 52322 194751 52325
rect 163700 52320 194751 52322
rect 163700 52264 194690 52320
rect 194746 52264 194751 52320
rect 163700 52262 194751 52264
rect 163700 52260 163706 52262
rect 194685 52259 194751 52262
rect 194685 51914 194751 51917
rect 405733 51914 405799 51917
rect 194685 51912 405799 51914
rect 194685 51856 194690 51912
rect 194746 51856 405738 51912
rect 405794 51856 405799 51912
rect 194685 51854 405799 51856
rect 194685 51851 194751 51854
rect 405733 51851 405799 51854
rect 27705 51778 27771 51781
rect 100753 51778 100819 51781
rect 27705 51776 100819 51778
rect 27705 51720 27710 51776
rect 27766 51720 100758 51776
rect 100814 51720 100819 51776
rect 27705 51718 100819 51720
rect 27705 51715 27771 51718
rect 100753 51715 100819 51718
rect 202781 51778 202847 51781
rect 455413 51778 455479 51781
rect 202781 51776 455479 51778
rect 202781 51720 202786 51776
rect 202842 51720 455418 51776
rect 455474 51720 455479 51776
rect 202781 51718 455479 51720
rect 202781 51715 202847 51718
rect 455413 51715 455479 51718
rect 100845 50962 100911 50965
rect 101857 50962 101923 50965
rect 134006 50962 134012 50964
rect 100845 50960 134012 50962
rect 100845 50904 100850 50960
rect 100906 50904 101862 50960
rect 101918 50904 134012 50960
rect 100845 50902 134012 50904
rect 100845 50899 100911 50902
rect 101857 50899 101923 50902
rect 134006 50900 134012 50902
rect 134076 50900 134082 50964
rect 165470 50900 165476 50964
rect 165540 50962 165546 50964
rect 198733 50962 198799 50965
rect 199561 50962 199627 50965
rect 203057 50964 203123 50965
rect 203006 50962 203012 50964
rect 165540 50960 199627 50962
rect 165540 50904 198738 50960
rect 198794 50904 199566 50960
rect 199622 50904 199627 50960
rect 165540 50902 199627 50904
rect 202966 50902 203012 50962
rect 203076 50960 203123 50964
rect 203118 50904 203123 50960
rect 165540 50900 165546 50902
rect 198733 50899 198799 50902
rect 199561 50899 199627 50902
rect 203006 50900 203012 50902
rect 203076 50900 203123 50904
rect 203057 50899 203123 50900
rect 158294 50764 158300 50828
rect 158364 50826 158370 50828
rect 190453 50826 190519 50829
rect 158364 50824 190519 50826
rect 158364 50768 190458 50824
rect 190514 50768 190519 50824
rect 158364 50766 190519 50768
rect 158364 50764 158370 50766
rect 190410 50763 190519 50766
rect 144678 50628 144684 50692
rect 144748 50690 144754 50692
rect 149789 50690 149855 50693
rect 144748 50688 149855 50690
rect 144748 50632 149794 50688
rect 149850 50632 149855 50688
rect 144748 50630 149855 50632
rect 144748 50628 144754 50630
rect 149789 50627 149855 50630
rect 190410 50418 190470 50763
rect 338113 50418 338179 50421
rect 190410 50416 338179 50418
rect 190410 50360 338118 50416
rect 338174 50360 338179 50416
rect 190410 50358 338179 50360
rect 338113 50355 338179 50358
rect 30373 50282 30439 50285
rect 100845 50282 100911 50285
rect 30373 50280 100911 50282
rect 30373 50224 30378 50280
rect 30434 50224 100850 50280
rect 100906 50224 100911 50280
rect 30373 50222 100911 50224
rect 30373 50219 30439 50222
rect 100845 50219 100911 50222
rect 199561 50282 199627 50285
rect 418797 50282 418863 50285
rect 199561 50280 418863 50282
rect 199561 50224 199566 50280
rect 199622 50224 418802 50280
rect 418858 50224 418863 50280
rect 199561 50222 418863 50224
rect 199561 50219 199627 50222
rect 418797 50219 418863 50222
rect 100845 49602 100911 49605
rect 101765 49602 101831 49605
rect 135478 49602 135484 49604
rect 100845 49600 135484 49602
rect 100845 49544 100850 49600
rect 100906 49544 101770 49600
rect 101826 49544 135484 49600
rect 100845 49542 135484 49544
rect 100845 49539 100911 49542
rect 101765 49539 101831 49542
rect 135478 49540 135484 49542
rect 135548 49540 135554 49604
rect 166574 49540 166580 49604
rect 166644 49602 166650 49604
rect 200113 49602 200179 49605
rect 201401 49602 201467 49605
rect 166644 49600 201467 49602
rect 166644 49544 200118 49600
rect 200174 49544 201406 49600
rect 201462 49544 201467 49600
rect 166644 49542 201467 49544
rect 166644 49540 166650 49542
rect 200113 49539 200179 49542
rect 201401 49539 201467 49542
rect 162710 49404 162716 49468
rect 162780 49466 162786 49468
rect 195973 49466 196039 49469
rect 162780 49464 196039 49466
rect 162780 49408 195978 49464
rect 196034 49408 196039 49464
rect 162780 49406 196039 49408
rect 162780 49404 162786 49406
rect 195973 49403 196039 49406
rect 159030 49268 159036 49332
rect 159100 49330 159106 49332
rect 159100 49270 200130 49330
rect 159100 49268 159106 49270
rect 190494 48996 190500 49060
rect 190564 49058 190570 49060
rect 190686 49058 190746 49270
rect 200070 49194 200130 49270
rect 356053 49194 356119 49197
rect 200070 49192 356119 49194
rect 200070 49136 356058 49192
rect 356114 49136 356119 49192
rect 200070 49134 356119 49136
rect 356053 49131 356119 49134
rect 190564 48998 190746 49058
rect 195973 49058 196039 49061
rect 387793 49058 387859 49061
rect 195973 49056 387859 49058
rect 195973 49000 195978 49056
rect 196034 49000 387798 49056
rect 387854 49000 387859 49056
rect 195973 48998 387859 49000
rect 190564 48996 190570 48998
rect 195973 48995 196039 48998
rect 387793 48995 387859 48998
rect 39297 48922 39363 48925
rect 100845 48922 100911 48925
rect 39297 48920 100911 48922
rect 39297 48864 39302 48920
rect 39358 48864 100850 48920
rect 100906 48864 100911 48920
rect 39297 48862 100911 48864
rect 39297 48859 39363 48862
rect 100845 48859 100911 48862
rect 201401 48922 201467 48925
rect 440233 48922 440299 48925
rect 201401 48920 440299 48922
rect 201401 48864 201406 48920
rect 201462 48864 440238 48920
rect 440294 48864 440299 48920
rect 201401 48862 440299 48864
rect 201401 48859 201467 48862
rect 440233 48859 440299 48862
rect 100845 48242 100911 48245
rect 101949 48242 102015 48245
rect 135846 48242 135852 48244
rect 100845 48240 135852 48242
rect 100845 48184 100850 48240
rect 100906 48184 101954 48240
rect 102010 48184 135852 48240
rect 100845 48182 135852 48184
rect 100845 48179 100911 48182
rect 101949 48179 102015 48182
rect 135846 48180 135852 48182
rect 135916 48180 135922 48244
rect 169334 48180 169340 48244
rect 169404 48242 169410 48244
rect 203333 48242 203399 48245
rect 204161 48242 204227 48245
rect 169404 48240 204227 48242
rect 169404 48184 203338 48240
rect 203394 48184 204166 48240
rect 204222 48184 204227 48240
rect 169404 48182 204227 48184
rect 169404 48180 169410 48182
rect 203333 48179 203399 48182
rect 204161 48179 204227 48182
rect 161238 48044 161244 48108
rect 161308 48106 161314 48108
rect 161308 48046 180810 48106
rect 161308 48044 161314 48046
rect 180750 47698 180810 48046
rect 194593 47698 194659 47701
rect 373993 47698 374059 47701
rect 180750 47696 374059 47698
rect 180750 47640 194598 47696
rect 194654 47640 373998 47696
rect 374054 47640 374059 47696
rect 180750 47638 374059 47640
rect 194593 47635 194659 47638
rect 373993 47635 374059 47638
rect 44173 47562 44239 47565
rect 100845 47562 100911 47565
rect 44173 47560 100911 47562
rect 44173 47504 44178 47560
rect 44234 47504 100850 47560
rect 100906 47504 100911 47560
rect 44173 47502 100911 47504
rect 44173 47499 44239 47502
rect 100845 47499 100911 47502
rect 204161 47562 204227 47565
rect 470593 47562 470659 47565
rect 204161 47560 470659 47562
rect 204161 47504 204166 47560
rect 204222 47504 470598 47560
rect 470654 47504 470659 47560
rect 204161 47502 470659 47504
rect 204161 47499 204227 47502
rect 470593 47499 470659 47502
rect 110505 46882 110571 46885
rect 110873 46882 110939 46885
rect 137686 46882 137692 46884
rect 110505 46880 137692 46882
rect 110505 46824 110510 46880
rect 110566 46824 110878 46880
rect 110934 46824 137692 46880
rect 110505 46822 137692 46824
rect 110505 46819 110571 46822
rect 110873 46819 110939 46822
rect 137686 46820 137692 46822
rect 137756 46820 137762 46884
rect 168046 46820 168052 46884
rect 168116 46882 168122 46884
rect 168116 46822 200130 46882
rect 168116 46820 168122 46822
rect 56593 46202 56659 46205
rect 110505 46202 110571 46205
rect 56593 46200 110571 46202
rect 56593 46144 56598 46200
rect 56654 46144 110510 46200
rect 110566 46144 110571 46200
rect 56593 46142 110571 46144
rect 200070 46202 200130 46822
rect 583520 46338 584960 46428
rect 583342 46278 584960 46338
rect 201534 46202 201540 46204
rect 200070 46142 201540 46202
rect 56593 46139 56659 46142
rect 110505 46139 110571 46142
rect 201534 46140 201540 46142
rect 201604 46202 201610 46204
rect 458173 46202 458239 46205
rect 201604 46200 458239 46202
rect 201604 46144 458178 46200
rect 458234 46144 458239 46200
rect 201604 46142 458239 46144
rect 583342 46202 583402 46278
rect 583520 46202 584960 46278
rect 583342 46188 584960 46202
rect 583342 46142 583586 46188
rect 201604 46140 201610 46142
rect 458173 46139 458239 46142
rect 142061 45660 142127 45661
rect 142061 45658 142108 45660
rect 142016 45656 142108 45658
rect 142172 45658 142178 45660
rect -960 45522 480 45612
rect 142016 45600 142066 45656
rect 142016 45598 142108 45600
rect 142061 45596 142108 45598
rect 142172 45598 142254 45658
rect 142172 45596 142178 45598
rect 192334 45596 192340 45660
rect 192404 45658 192410 45660
rect 583526 45658 583586 46142
rect 192404 45598 583586 45658
rect 192404 45596 192410 45598
rect 142061 45595 142127 45596
rect 3417 45522 3483 45525
rect 142061 45524 142127 45525
rect 142061 45522 142108 45524
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect 142016 45520 142108 45522
rect 142172 45522 142178 45524
rect 142016 45464 142066 45520
rect 142016 45462 142108 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 142061 45460 142108 45462
rect 142172 45462 142254 45522
rect 142172 45460 142178 45462
rect 142061 45459 142127 45460
rect 146702 44916 146708 44980
rect 146772 44978 146778 44980
rect 194593 44978 194659 44981
rect 146772 44976 194659 44978
rect 146772 44920 194598 44976
rect 194654 44920 194659 44976
rect 146772 44918 194659 44920
rect 146772 44916 146778 44918
rect 194593 44915 194659 44918
rect 151118 44780 151124 44844
rect 151188 44842 151194 44844
rect 249793 44842 249859 44845
rect 151188 44840 249859 44842
rect 151188 44784 249798 44840
rect 249854 44784 249859 44840
rect 151188 44782 249859 44784
rect 151188 44780 151194 44782
rect 249793 44779 249859 44782
rect 108389 44162 108455 44165
rect 138054 44162 138060 44164
rect 108389 44160 138060 44162
rect 108389 44104 108394 44160
rect 108450 44104 138060 44160
rect 108389 44102 138060 44104
rect 108389 44099 108455 44102
rect 138054 44100 138060 44102
rect 138124 44100 138130 44164
rect 166758 44100 166764 44164
rect 166828 44162 166834 44164
rect 200665 44162 200731 44165
rect 166828 44160 209790 44162
rect 166828 44104 200670 44160
rect 200726 44104 209790 44160
rect 166828 44102 209790 44104
rect 166828 44100 166834 44102
rect 200665 44099 200731 44102
rect 169518 43964 169524 44028
rect 169588 44026 169594 44028
rect 202873 44026 202939 44029
rect 169588 44024 202939 44026
rect 169588 43968 202878 44024
rect 202934 43968 202939 44024
rect 169588 43966 202939 43968
rect 169588 43964 169594 43966
rect 202873 43963 202939 43966
rect 209730 43618 209790 44102
rect 427813 43618 427879 43621
rect 209730 43616 427879 43618
rect 209730 43560 427818 43616
rect 427874 43560 427879 43616
rect 209730 43558 427879 43560
rect 427813 43555 427879 43558
rect 74533 43482 74599 43485
rect 108389 43482 108455 43485
rect 74533 43480 108455 43482
rect 74533 43424 74538 43480
rect 74594 43424 108394 43480
rect 108450 43424 108455 43480
rect 74533 43422 108455 43424
rect 74533 43419 74599 43422
rect 108389 43419 108455 43422
rect 202873 43482 202939 43485
rect 476113 43482 476179 43485
rect 202873 43480 476179 43482
rect 202873 43424 202878 43480
rect 202934 43424 476118 43480
rect 476174 43424 476179 43480
rect 202873 43422 476179 43424
rect 202873 43419 202939 43422
rect 476113 43419 476179 43422
rect 149278 42060 149284 42124
rect 149348 42122 149354 42124
rect 230473 42122 230539 42125
rect 149348 42120 230539 42122
rect 149348 42064 230478 42120
rect 230534 42064 230539 42120
rect 149348 42062 230539 42064
rect 149348 42060 149354 42062
rect 230473 42059 230539 42062
rect 152958 40564 152964 40628
rect 153028 40626 153034 40628
rect 267733 40626 267799 40629
rect 153028 40624 267799 40626
rect 153028 40568 267738 40624
rect 267794 40568 267799 40624
rect 153028 40566 267799 40568
rect 153028 40564 153034 40566
rect 267733 40563 267799 40566
rect 17309 36546 17375 36549
rect 133454 36546 133460 36548
rect 17309 36544 133460 36546
rect 17309 36488 17314 36544
rect 17370 36488 133460 36544
rect 17309 36486 133460 36488
rect 17309 36483 17375 36486
rect 133454 36484 133460 36486
rect 133524 36484 133530 36548
rect 170990 36484 170996 36548
rect 171060 36546 171066 36548
rect 494053 36546 494119 36549
rect 171060 36544 494119 36546
rect 171060 36488 494058 36544
rect 494114 36488 494119 36544
rect 171060 36486 494119 36488
rect 171060 36484 171066 36486
rect 494053 36483 494119 36486
rect 142102 36076 142108 36140
rect 142172 36076 142178 36140
rect 142110 36005 142170 36076
rect 142061 36002 142170 36005
rect 142016 36000 142170 36002
rect 142016 35944 142066 36000
rect 142122 35944 142170 36000
rect 142016 35942 142170 35944
rect 142061 35939 142127 35942
rect 142061 35866 142127 35869
rect 142286 35866 142292 35868
rect 142016 35864 142292 35866
rect 142016 35808 142066 35864
rect 142122 35808 142292 35864
rect 142016 35806 142292 35808
rect 142061 35803 142127 35806
rect 142286 35804 142292 35806
rect 142356 35804 142362 35868
rect 24853 33826 24919 33829
rect 134926 33826 134932 33828
rect 24853 33824 134932 33826
rect 24853 33768 24858 33824
rect 24914 33768 134932 33824
rect 24853 33766 134932 33768
rect 24853 33763 24919 33766
rect 134926 33764 134932 33766
rect 134996 33764 135002 33828
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect -960 32406 674 32466
rect -960 32330 480 32406
rect 614 32330 674 32406
rect 148910 32404 148916 32468
rect 148980 32466 148986 32468
rect 212533 32466 212599 32469
rect 148980 32464 212599 32466
rect 148980 32408 212538 32464
rect 212594 32408 212599 32464
rect 148980 32406 212599 32408
rect 148980 32404 148986 32406
rect 212533 32403 212599 32406
rect -960 32316 674 32330
rect 246 32270 674 32316
rect 246 31786 306 32270
rect 120574 31786 120580 31788
rect 246 31726 120580 31786
rect 120574 31724 120580 31726
rect 120644 31724 120650 31788
rect 145414 26964 145420 27028
rect 145484 27026 145490 27028
rect 171777 27026 171843 27029
rect 145484 27024 171843 27026
rect 145484 26968 171782 27024
rect 171838 26968 171843 27024
rect 145484 26966 171843 26968
rect 145484 26964 145490 26966
rect 171777 26963 171843 26966
rect 152406 26828 152412 26892
rect 152476 26890 152482 26892
rect 264973 26890 265039 26893
rect 152476 26888 265039 26890
rect 152476 26832 264978 26888
rect 265034 26832 265039 26888
rect 152476 26830 265039 26832
rect 152476 26828 152482 26830
rect 264973 26827 265039 26830
rect 142061 26348 142127 26349
rect 142061 26346 142108 26348
rect 142016 26344 142108 26346
rect 142172 26346 142178 26348
rect 142016 26288 142066 26344
rect 142016 26286 142108 26288
rect 142061 26284 142108 26286
rect 142172 26286 142254 26346
rect 142172 26284 142178 26286
rect 142061 26283 142127 26284
rect 142061 26212 142127 26213
rect 142061 26210 142108 26212
rect 142016 26208 142108 26210
rect 142172 26210 142178 26212
rect 142016 26152 142066 26208
rect 142016 26150 142108 26152
rect 142061 26148 142108 26150
rect 142172 26150 142254 26210
rect 142172 26148 142178 26150
rect 142061 26147 142127 26148
rect 144494 21252 144500 21316
rect 144564 21314 144570 21316
rect 158713 21314 158779 21317
rect 144564 21312 158779 21314
rect 144564 21256 158718 21312
rect 158774 21256 158779 21312
rect 144564 21254 158779 21256
rect 144564 21252 144570 21254
rect 158713 21251 158779 21254
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 116526 19410 116532 19412
rect -960 19350 116532 19410
rect -960 19260 480 19350
rect 116526 19348 116532 19350
rect 116596 19348 116602 19412
rect 149646 18532 149652 18596
rect 149716 18594 149722 18596
rect 229093 18594 229159 18597
rect 149716 18592 229159 18594
rect 149716 18536 229098 18592
rect 229154 18536 229159 18592
rect 149716 18534 229159 18536
rect 149716 18532 149722 18534
rect 229093 18531 229159 18534
rect 142061 16690 142127 16693
rect 142286 16690 142292 16692
rect 142016 16688 142292 16690
rect 142016 16632 142066 16688
rect 142122 16632 142292 16688
rect 142016 16630 142292 16632
rect 142061 16627 142127 16630
rect 142286 16628 142292 16630
rect 142356 16628 142362 16692
rect 142061 16554 142127 16557
rect 142016 16552 142170 16554
rect 142016 16496 142066 16552
rect 142122 16496 142170 16552
rect 142016 16494 142170 16496
rect 142061 16491 142170 16494
rect 142110 16420 142170 16491
rect 142102 16356 142108 16420
rect 142172 16356 142178 16420
rect 144310 15812 144316 15876
rect 144380 15874 144386 15876
rect 160093 15874 160159 15877
rect 144380 15872 160159 15874
rect 144380 15816 160098 15872
rect 160154 15816 160159 15872
rect 144380 15814 160159 15816
rect 144380 15812 144386 15814
rect 160093 15811 160159 15814
rect 158478 11596 158484 11660
rect 158548 11658 158554 11660
rect 336273 11658 336339 11661
rect 158548 11656 336339 11658
rect 158548 11600 336278 11656
rect 336334 11600 336339 11656
rect 158548 11598 336339 11600
rect 158548 11596 158554 11598
rect 336273 11595 336339 11598
rect 142061 7036 142127 7037
rect 142061 7034 142108 7036
rect 142016 7032 142108 7034
rect 142172 7034 142178 7036
rect 142016 6976 142066 7032
rect 142016 6974 142108 6976
rect 142061 6972 142108 6974
rect 142172 6974 142254 7034
rect 142172 6972 142178 6974
rect 142061 6971 142127 6972
rect 142061 6900 142127 6901
rect 142061 6898 142108 6900
rect 142016 6896 142108 6898
rect 142172 6898 142178 6900
rect 142016 6840 142066 6896
rect 142016 6838 142108 6840
rect 142061 6836 142108 6838
rect 142172 6838 142254 6898
rect 142172 6836 142178 6838
rect 142061 6835 142127 6836
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 144126 4796 144132 4860
rect 144196 4858 144202 4860
rect 161289 4858 161355 4861
rect 144196 4856 161355 4858
rect 144196 4800 161294 4856
rect 161350 4800 161355 4856
rect 144196 4798 161355 4800
rect 144196 4796 144202 4798
rect 161289 4795 161355 4798
rect 111609 3362 111675 3365
rect 142061 3362 142127 3365
rect 111609 3360 142127 3362
rect 111609 3304 111614 3360
rect 111670 3304 142066 3360
rect 142122 3304 142127 3360
rect 111609 3302 142127 3304
rect 111609 3299 111675 3302
rect 142061 3299 142127 3302
<< via3 >>
rect 189028 278020 189092 278084
rect 189028 277476 189092 277540
rect 189212 275980 189276 276044
rect 197492 265372 197556 265436
rect 196204 265236 196268 265300
rect 111564 265100 111628 265164
rect 113036 264964 113100 265028
rect 194548 265100 194612 265164
rect 197676 264964 197740 265028
rect 119844 263876 119908 263940
rect 121316 263740 121380 263804
rect 112852 263604 112916 263668
rect 114140 262924 114204 262988
rect 115612 262788 115676 262852
rect 112668 262652 112732 262716
rect 113956 262516 114020 262580
rect 116716 262380 116780 262444
rect 193444 262652 193508 262716
rect 191972 262516 192036 262580
rect 193628 262380 193692 262444
rect 115428 262244 115492 262308
rect 190500 262244 190564 262308
rect 192156 262244 192220 262308
rect 111380 261020 111444 261084
rect 111196 260884 111260 260948
rect 117084 260340 117148 260404
rect 121132 260204 121196 260268
rect 118372 260068 118436 260132
rect 116900 259932 116964 259996
rect 189580 260068 189644 260132
rect 118188 259796 118252 259860
rect 113772 259660 113836 259724
rect 191788 259660 191852 259724
rect 115796 259524 115860 259588
rect 186084 259524 186148 259588
rect 186084 212468 186148 212532
rect 187188 212468 187252 212532
rect 141556 200636 141620 200700
rect 136588 200500 136652 200564
rect 138060 200364 138124 200428
rect 150204 200228 150268 200292
rect 170260 200228 170324 200292
rect 133644 200092 133708 200156
rect 138060 200092 138124 200156
rect 138612 199956 138676 200020
rect 133092 199820 133156 199884
rect 133644 199880 133708 199884
rect 133644 199824 133648 199880
rect 133648 199824 133704 199880
rect 133704 199824 133708 199880
rect 133644 199820 133708 199824
rect 134748 199820 134812 199884
rect 136036 199820 136100 199884
rect 136404 199684 136468 199748
rect 137140 199684 137204 199748
rect 138796 199820 138860 199884
rect 137692 199684 137756 199748
rect 140636 199820 140700 199884
rect 141004 199880 141068 199884
rect 141004 199824 141008 199880
rect 141008 199824 141064 199880
rect 141064 199824 141068 199880
rect 141004 199820 141068 199824
rect 142476 199858 142480 199884
rect 142480 199858 142536 199884
rect 142536 199858 142540 199884
rect 142476 199820 142540 199858
rect 144500 199858 144504 199884
rect 144504 199858 144560 199884
rect 144560 199858 144564 199884
rect 144500 199820 144564 199858
rect 145420 199858 145424 199884
rect 145424 199858 145480 199884
rect 145480 199858 145484 199884
rect 145420 199820 145484 199858
rect 147076 199820 147140 199884
rect 147812 199880 147876 199884
rect 147812 199824 147816 199880
rect 147816 199824 147872 199880
rect 147872 199824 147876 199880
rect 147812 199820 147876 199824
rect 147996 199858 148000 199884
rect 148000 199858 148056 199884
rect 148056 199858 148060 199884
rect 147996 199820 148060 199858
rect 148548 199820 148612 199884
rect 140084 199684 140148 199748
rect 140820 199744 140884 199748
rect 140820 199688 140824 199744
rect 140824 199688 140880 199744
rect 140880 199688 140884 199744
rect 140820 199684 140884 199688
rect 145604 199684 145668 199748
rect 136588 199608 136652 199612
rect 136588 199552 136638 199608
rect 136638 199552 136652 199608
rect 136588 199548 136652 199552
rect 139348 199548 139412 199612
rect 141556 199548 141620 199612
rect 148732 199744 148796 199748
rect 150020 200092 150084 200156
rect 149652 199858 149656 199884
rect 149656 199858 149712 199884
rect 149712 199858 149716 199884
rect 149652 199820 149716 199858
rect 150388 199820 150452 199884
rect 150756 199858 150760 199884
rect 150760 199858 150816 199884
rect 150816 199858 150820 199884
rect 151308 199956 151372 200020
rect 151492 199956 151556 200020
rect 153516 199956 153580 200020
rect 150756 199820 150820 199858
rect 152044 199880 152108 199884
rect 152044 199824 152048 199880
rect 152048 199824 152104 199880
rect 152104 199824 152108 199880
rect 152044 199820 152108 199824
rect 152228 199820 152292 199884
rect 152780 199858 152784 199884
rect 152784 199858 152840 199884
rect 152840 199858 152844 199884
rect 152780 199820 152844 199858
rect 153148 199820 153212 199884
rect 153332 199820 153396 199884
rect 153884 199820 153948 199884
rect 154804 199880 154868 199884
rect 154804 199824 154808 199880
rect 154808 199824 154864 199880
rect 154864 199824 154868 199880
rect 154804 199820 154868 199824
rect 155540 199820 155604 199884
rect 156092 199820 156156 199884
rect 157380 199820 157444 199884
rect 165292 199956 165356 200020
rect 160508 199820 160572 199884
rect 162348 199820 162412 199884
rect 163452 199880 163516 199884
rect 163452 199824 163456 199880
rect 163456 199824 163512 199880
rect 163512 199824 163516 199880
rect 163452 199820 163516 199824
rect 163636 199820 163700 199884
rect 164372 199820 164436 199884
rect 165108 199880 165172 199884
rect 165108 199824 165112 199880
rect 165112 199824 165168 199880
rect 165168 199824 165172 199880
rect 165108 199820 165172 199824
rect 168788 199956 168852 200020
rect 174676 199956 174740 200020
rect 166580 199820 166644 199884
rect 167132 199880 167196 199884
rect 167132 199824 167136 199880
rect 167136 199824 167192 199880
rect 167192 199824 167196 199880
rect 167132 199820 167196 199824
rect 167546 199820 167610 199884
rect 167868 199880 167932 199884
rect 167868 199824 167872 199880
rect 167872 199824 167928 199880
rect 167928 199824 167932 199880
rect 167868 199820 167932 199824
rect 168972 199820 169036 199884
rect 170812 199820 170876 199884
rect 171364 199820 171428 199884
rect 171548 199880 171612 199884
rect 171548 199824 171552 199880
rect 171552 199824 171608 199880
rect 171608 199824 171612 199880
rect 171548 199820 171612 199824
rect 172468 199880 172532 199884
rect 172468 199824 172472 199880
rect 172472 199824 172528 199880
rect 172528 199824 172532 199880
rect 172468 199820 172532 199824
rect 172652 199820 172716 199884
rect 174492 199820 174556 199884
rect 175044 199880 175108 199884
rect 175044 199824 175048 199880
rect 175048 199824 175104 199880
rect 175104 199824 175108 199880
rect 175044 199820 175108 199824
rect 175596 199880 175660 199884
rect 175596 199824 175600 199880
rect 175600 199824 175656 199880
rect 175656 199824 175660 199880
rect 175596 199820 175660 199824
rect 176332 199820 176396 199884
rect 148732 199688 148736 199744
rect 148736 199688 148792 199744
rect 148792 199688 148796 199744
rect 148732 199684 148796 199688
rect 182772 199684 182836 199748
rect 180748 199548 180812 199612
rect 122604 199412 122668 199476
rect 149652 199472 149716 199476
rect 149652 199416 149666 199472
rect 149666 199416 149716 199472
rect 149652 199412 149716 199416
rect 150204 199412 150268 199476
rect 151676 199472 151740 199476
rect 151676 199416 151726 199472
rect 151726 199416 151740 199472
rect 151676 199412 151740 199416
rect 152044 199412 152108 199476
rect 156828 199412 156892 199476
rect 153884 199276 153948 199340
rect 154804 199276 154868 199340
rect 156092 199276 156156 199340
rect 157380 199276 157444 199340
rect 158300 199276 158364 199340
rect 161244 199276 161308 199340
rect 165108 199336 165172 199340
rect 165108 199280 165158 199336
rect 165158 199280 165172 199336
rect 165108 199276 165172 199280
rect 170260 199276 170324 199340
rect 170444 199336 170508 199340
rect 170444 199280 170458 199336
rect 170458 199280 170508 199336
rect 170444 199276 170508 199280
rect 170812 199336 170876 199340
rect 170812 199280 170862 199336
rect 170862 199280 170876 199336
rect 170812 199276 170876 199280
rect 171364 199276 171428 199340
rect 171732 199276 171796 199340
rect 174492 199412 174556 199476
rect 174676 199412 174740 199476
rect 175596 199412 175660 199476
rect 176516 199412 176580 199476
rect 179644 199140 179708 199204
rect 135852 199004 135916 199068
rect 136404 199064 136468 199068
rect 136404 199008 136454 199064
rect 136454 199008 136468 199064
rect 136404 199004 136468 199008
rect 139348 199064 139412 199068
rect 139348 199008 139362 199064
rect 139362 199008 139412 199064
rect 139348 199004 139412 199008
rect 140268 199004 140332 199068
rect 145420 199004 145484 199068
rect 146892 198868 146956 198932
rect 147996 198928 148060 198932
rect 147996 198872 148010 198928
rect 148010 198872 148060 198928
rect 147996 198868 148060 198872
rect 148732 198868 148796 198932
rect 157196 198868 157260 198932
rect 139164 198732 139228 198796
rect 150756 198732 150820 198796
rect 157012 198792 157076 198796
rect 157012 198736 157026 198792
rect 157026 198736 157076 198792
rect 157012 198732 157076 198736
rect 158116 198732 158180 198796
rect 166396 199004 166460 199068
rect 175964 199004 176028 199068
rect 176516 199064 176580 199068
rect 176516 199008 176530 199064
rect 176530 199008 176580 199064
rect 176516 199004 176580 199008
rect 166028 198928 166092 198932
rect 166028 198872 166042 198928
rect 166042 198872 166092 198928
rect 166028 198868 166092 198872
rect 166212 198868 166276 198932
rect 167868 198928 167932 198932
rect 167868 198872 167882 198928
rect 167882 198872 167932 198928
rect 167868 198868 167932 198872
rect 178356 198868 178420 198932
rect 172468 198732 172532 198796
rect 199332 198732 199396 198796
rect 133460 198656 133524 198660
rect 133460 198600 133510 198656
rect 133510 198600 133524 198656
rect 133460 198596 133524 198600
rect 130884 198460 130948 198524
rect 148916 198596 148980 198660
rect 150388 198460 150452 198524
rect 125364 198324 125428 198388
rect 125180 198188 125244 198252
rect 124996 198052 125060 198116
rect 134380 197976 134444 197980
rect 134380 197920 134430 197976
rect 134430 197920 134444 197976
rect 134380 197916 134444 197920
rect 134564 197916 134628 197980
rect 137508 197916 137572 197980
rect 133644 197780 133708 197844
rect 134932 197780 134996 197844
rect 136588 197780 136652 197844
rect 145604 198188 145668 198252
rect 157564 198188 157628 198252
rect 139348 198112 139412 198116
rect 139348 198056 139398 198112
rect 139398 198056 139412 198112
rect 139348 198052 139412 198056
rect 140084 198052 140148 198116
rect 140452 198052 140516 198116
rect 144132 198052 144196 198116
rect 166580 198112 166644 198116
rect 187004 198596 187068 198660
rect 175596 198460 175660 198524
rect 187740 198460 187804 198524
rect 169892 198188 169956 198252
rect 189396 198324 189460 198388
rect 198964 198188 199028 198252
rect 166580 198056 166594 198112
rect 166594 198056 166644 198112
rect 166580 198052 166644 198056
rect 176700 198052 176764 198116
rect 177068 198052 177132 198116
rect 141004 197916 141068 197980
rect 142660 197916 142724 197980
rect 144684 197916 144748 197980
rect 133276 197704 133340 197708
rect 133276 197648 133326 197704
rect 133326 197648 133340 197704
rect 133276 197644 133340 197648
rect 160508 197644 160572 197708
rect 169156 197916 169220 197980
rect 174124 197916 174188 197980
rect 174492 197916 174556 197980
rect 176884 197916 176948 197980
rect 187924 197780 187988 197844
rect 179460 197644 179524 197708
rect 130700 197508 130764 197572
rect 148732 197508 148796 197572
rect 162164 197508 162228 197572
rect 164556 197508 164620 197572
rect 167684 197508 167748 197572
rect 174860 197508 174924 197572
rect 176700 197508 176764 197572
rect 180932 197508 180996 197572
rect 126652 197432 126716 197436
rect 126652 197376 126702 197432
rect 126702 197376 126716 197432
rect 126652 197372 126716 197376
rect 130516 197372 130580 197436
rect 153332 197372 153396 197436
rect 126836 197236 126900 197300
rect 156644 197236 156708 197300
rect 157196 197372 157260 197436
rect 160876 197372 160940 197436
rect 163084 197372 163148 197436
rect 164924 197372 164988 197436
rect 168052 197432 168116 197436
rect 168052 197376 168066 197432
rect 168066 197376 168116 197432
rect 168052 197372 168116 197376
rect 169524 197372 169588 197436
rect 170076 197372 170140 197436
rect 171364 197372 171428 197436
rect 171916 197372 171980 197436
rect 172836 197372 172900 197436
rect 174308 197372 174372 197436
rect 175412 197372 175476 197436
rect 161060 197296 161124 197300
rect 161060 197240 161074 197296
rect 161074 197240 161124 197296
rect 161060 197236 161124 197240
rect 163268 197236 163332 197300
rect 165108 197236 165172 197300
rect 165292 197296 165356 197300
rect 165292 197240 165342 197296
rect 165342 197240 165356 197296
rect 165292 197236 165356 197240
rect 165660 197236 165724 197300
rect 167316 197236 167380 197300
rect 169340 197236 169404 197300
rect 170444 197296 170508 197300
rect 170444 197240 170458 197296
rect 170458 197240 170508 197296
rect 170444 197236 170508 197240
rect 173020 197296 173084 197300
rect 173020 197240 173034 197296
rect 173034 197240 173084 197296
rect 173020 197236 173084 197240
rect 173388 197236 173452 197300
rect 175044 197296 175108 197300
rect 175044 197240 175058 197296
rect 175058 197240 175108 197296
rect 175044 197236 175108 197240
rect 175780 197236 175844 197300
rect 160508 197100 160572 197164
rect 193260 197100 193324 197164
rect 140820 196964 140884 197028
rect 143580 196964 143644 197028
rect 149836 196964 149900 197028
rect 151308 196964 151372 197028
rect 178172 196964 178236 197028
rect 149468 196828 149532 196892
rect 151676 196692 151740 196756
rect 157932 196692 157996 196756
rect 158852 196692 158916 196756
rect 161980 196692 162044 196756
rect 118556 196556 118620 196620
rect 159036 196556 159100 196620
rect 168788 196556 168852 196620
rect 142476 196420 142540 196484
rect 149652 196420 149716 196484
rect 133092 196148 133156 196212
rect 131620 196012 131684 196076
rect 133276 196012 133340 196076
rect 140820 196012 140884 196076
rect 145236 196012 145300 196076
rect 147812 196012 147876 196076
rect 151492 196012 151556 196076
rect 131804 195876 131868 195940
rect 148548 195876 148612 195940
rect 198780 195876 198844 195940
rect 128124 195740 128188 195804
rect 197308 195740 197372 195804
rect 132172 195604 132236 195668
rect 151124 195604 151188 195668
rect 156276 195604 156340 195668
rect 200620 195604 200684 195668
rect 126468 195468 126532 195532
rect 147260 195468 147324 195532
rect 176332 195468 176396 195532
rect 200988 195468 201052 195532
rect 142844 195332 142908 195396
rect 144684 195332 144748 195396
rect 182588 195332 182652 195396
rect 124076 195196 124140 195260
rect 200804 195196 200868 195260
rect 196020 195060 196084 195124
rect 124812 194108 124876 194172
rect 130332 193972 130396 194036
rect 155724 193972 155788 194036
rect 201724 193972 201788 194036
rect 201540 193836 201604 193900
rect 144500 193156 144564 193220
rect 167132 193156 167196 193220
rect 153700 191252 153764 191316
rect 136220 191116 136284 191180
rect 148180 191116 148244 191180
rect 163452 191116 163516 191180
rect 164372 191116 164436 191180
rect 164740 191176 164804 191180
rect 164740 191120 164754 191176
rect 164754 191120 164804 191176
rect 164740 191116 164804 191120
rect 135484 190980 135548 191044
rect 148364 190980 148428 191044
rect 154068 190844 154132 190908
rect 160508 190572 160572 190636
rect 161244 190572 161308 190636
rect 160692 190496 160756 190500
rect 160692 190440 160742 190496
rect 160742 190440 160756 190496
rect 160692 190436 160756 190440
rect 161428 190164 161492 190228
rect 143580 189620 143644 189684
rect 153884 189408 153948 189412
rect 153884 189352 153898 189408
rect 153898 189352 153948 189408
rect 153884 189348 153948 189352
rect 164004 189348 164068 189412
rect 141004 188804 141068 188868
rect 152412 183500 152476 183564
rect 138980 183228 139044 183292
rect 161428 180840 161492 180844
rect 161428 180784 161442 180840
rect 161442 180784 161492 180840
rect 161428 180780 161492 180784
rect 161428 180508 161492 180572
rect 161428 171184 161492 171188
rect 161428 171128 161442 171184
rect 161442 171128 161492 171184
rect 161428 171124 161492 171128
rect 161428 170852 161492 170916
rect 161428 161528 161492 161532
rect 161428 161472 161442 161528
rect 161442 161472 161492 161528
rect 161428 161468 161492 161472
rect 161428 161196 161492 161260
rect 186084 152628 186148 152692
rect 185164 152492 185228 152556
rect 185348 152356 185412 152420
rect 161428 151872 161492 151876
rect 161428 151816 161442 151872
rect 161442 151816 161492 151872
rect 161428 151812 161492 151816
rect 161428 151540 161492 151604
rect 203012 150316 203076 150380
rect 182956 150180 183020 150244
rect 181116 150044 181180 150108
rect 183140 149908 183204 149972
rect 183508 149772 183572 149836
rect 142476 149636 142540 149700
rect 184980 149636 185044 149700
rect 122420 147732 122484 147796
rect 201172 147732 201236 147796
rect 193812 147596 193876 147660
rect 196388 147460 196452 147524
rect 181300 147324 181364 147388
rect 198044 147188 198108 147252
rect 180012 147052 180076 147116
rect 183692 146916 183756 146980
rect 195100 146916 195164 146980
rect 115428 146236 115492 146300
rect 197860 146236 197924 146300
rect 111564 146100 111628 146164
rect 192524 146100 192588 146164
rect 111196 145964 111260 146028
rect 193996 145964 194060 146028
rect 113772 145828 113836 145892
rect 196572 145828 196636 145892
rect 114140 145692 114204 145756
rect 179828 145692 179892 145756
rect 113956 145556 114020 145620
rect 197676 145556 197740 145620
rect 120764 144876 120828 144940
rect 193628 144876 193692 144940
rect 118188 144740 118252 144804
rect 197492 144740 197556 144804
rect 144132 144604 144196 144668
rect 196204 144604 196268 144668
rect 112668 144468 112732 144532
rect 194548 144468 194612 144532
rect 112852 144332 112916 144396
rect 193444 144332 193508 144396
rect 118188 144196 118252 144260
rect 190500 144196 190564 144260
rect 116716 144060 116780 144124
rect 192156 144060 192220 144124
rect 115612 143924 115676 143988
rect 191972 143924 192036 143988
rect 113036 143788 113100 143852
rect 111380 143244 111444 143308
rect 187188 143380 187252 143444
rect 121132 143108 121196 143172
rect 121316 142972 121380 143036
rect 119844 142836 119908 142900
rect 189028 142836 189092 142900
rect 189580 142700 189644 142764
rect 189212 142564 189276 142628
rect 161612 142292 161676 142356
rect 122972 142156 123036 142220
rect 191788 142020 191852 142084
rect 117084 141748 117148 141812
rect 118372 141612 118436 141676
rect 116900 141476 116964 141540
rect 190500 141476 190564 141540
rect 115796 141340 115860 141404
rect 183876 141340 183940 141404
rect 141372 141204 141436 141268
rect 177804 141204 177868 141268
rect 141556 141068 141620 141132
rect 177436 141068 177500 141132
rect 188292 140932 188356 140996
rect 192340 140796 192404 140860
rect 190868 140720 190932 140724
rect 190868 140664 190882 140720
rect 190882 140664 190932 140720
rect 120580 140524 120644 140588
rect 190868 140660 190932 140664
rect 116532 140388 116596 140452
rect 184428 140448 184492 140452
rect 184428 140392 184442 140448
rect 184442 140392 184492 140448
rect 184428 140388 184492 140392
rect 191604 140252 191668 140316
rect 122236 140116 122300 140180
rect 188476 140116 188540 140180
rect 178908 139980 178972 140044
rect 119292 139844 119356 139908
rect 178540 139708 178604 139772
rect 189580 139844 189644 139908
rect 191972 139844 192036 139908
rect 185716 139768 185780 139772
rect 185716 139712 185766 139768
rect 185766 139712 185780 139768
rect 185716 139708 185780 139712
rect 189028 139708 189092 139772
rect 183324 139436 183388 139500
rect 122052 139300 122116 139364
rect 126284 139300 126348 139364
rect 127940 139300 128004 139364
rect 131988 139300 132052 139364
rect 150756 139300 150820 139364
rect 155356 139300 155420 139364
rect 154804 139164 154868 139228
rect 159220 139300 159284 139364
rect 159956 139300 160020 139364
rect 185716 139028 185780 139092
rect 183324 138892 183388 138956
rect 184428 138348 184492 138412
rect 186268 138212 186332 138276
rect 187188 138076 187252 138140
rect 122236 137940 122300 138004
rect 122788 137940 122852 138004
rect 185348 137940 185412 138004
rect 185164 137804 185228 137868
rect 122788 128420 122852 128484
rect 186084 127604 186148 127668
rect 188476 125564 188540 125628
rect 122788 123116 122852 123180
rect 122788 122436 122852 122500
rect 122788 113460 122852 113524
rect 122788 112780 122852 112844
rect 189580 111828 189644 111892
rect 122788 103804 122852 103868
rect 122788 103124 122852 103188
rect 122788 94148 122852 94212
rect 122788 93468 122852 93532
rect 122788 89660 122852 89724
rect 119292 84220 119356 84284
rect 134564 81908 134628 81972
rect 135116 81908 135180 81972
rect 139348 81500 139412 81564
rect 137324 81364 137388 81428
rect 142844 81364 142908 81428
rect 130700 81228 130764 81292
rect 143212 81228 143276 81292
rect 176516 81228 176580 81292
rect 130516 81092 130580 81156
rect 143396 81092 143460 81156
rect 173204 81092 173268 81156
rect 127940 80956 128004 81020
rect 147996 80956 148060 81020
rect 175228 80956 175292 81020
rect 124996 80820 125060 80884
rect 144868 80820 144932 80884
rect 160324 80820 160388 80884
rect 132172 80548 132236 80612
rect 170444 80684 170508 80748
rect 122788 80276 122852 80340
rect 126284 80276 126348 80340
rect 145052 80412 145116 80476
rect 138244 80276 138308 80340
rect 122972 80004 123036 80068
rect 134380 80004 134444 80068
rect 132908 79868 132972 79932
rect 145420 80004 145484 80068
rect 134564 79868 134628 79932
rect 131620 79732 131684 79796
rect 133092 79732 133156 79796
rect 133644 79732 133708 79796
rect 134748 79732 134812 79796
rect 135852 79868 135916 79932
rect 135116 79770 135120 79796
rect 135120 79770 135176 79796
rect 135176 79770 135180 79796
rect 135116 79732 135180 79770
rect 133276 79596 133340 79660
rect 134196 79596 134260 79660
rect 137140 79868 137204 79932
rect 137508 79868 137572 79932
rect 137692 79868 137756 79932
rect 136956 79732 137020 79796
rect 137324 79732 137388 79796
rect 134932 79596 134996 79660
rect 136220 79596 136284 79660
rect 136588 79596 136652 79660
rect 138980 79868 139044 79932
rect 139532 79928 139596 79932
rect 139532 79872 139536 79928
rect 139536 79872 139592 79928
rect 139592 79872 139596 79928
rect 139532 79868 139596 79872
rect 138796 79732 138860 79796
rect 139348 79732 139412 79796
rect 141004 79868 141068 79932
rect 138428 79596 138492 79660
rect 138612 79596 138676 79660
rect 139164 79656 139228 79660
rect 139164 79600 139214 79656
rect 139214 79600 139228 79656
rect 139164 79596 139228 79600
rect 139716 79656 139780 79660
rect 140268 79732 140332 79796
rect 143028 79868 143092 79932
rect 144316 79868 144380 79932
rect 145052 79868 145116 79932
rect 145420 79868 145484 79932
rect 164188 80548 164252 80612
rect 161244 80412 161308 80476
rect 176332 80548 176396 80612
rect 179644 80744 179708 80748
rect 179644 80688 179658 80744
rect 179658 80688 179708 80744
rect 179644 80684 179708 80688
rect 198964 80684 199028 80748
rect 156644 80276 156708 80340
rect 157196 80276 157260 80340
rect 160876 80276 160940 80340
rect 150756 80140 150820 80204
rect 154804 80140 154868 80204
rect 141004 79732 141068 79796
rect 141556 79732 141620 79796
rect 139716 79600 139730 79656
rect 139730 79600 139780 79656
rect 139716 79596 139780 79600
rect 140636 79596 140700 79660
rect 141372 79656 141436 79660
rect 141372 79600 141422 79656
rect 141422 79600 141436 79656
rect 141372 79596 141436 79600
rect 144500 79732 144564 79796
rect 144868 79732 144932 79796
rect 146892 79596 146956 79660
rect 148594 79906 148644 79932
rect 148644 79906 148658 79932
rect 148594 79868 148658 79906
rect 147996 79792 148060 79796
rect 147996 79736 148046 79792
rect 148046 79736 148060 79792
rect 147996 79732 148060 79736
rect 148364 79732 148428 79796
rect 149100 79732 149164 79796
rect 150204 79928 150268 79932
rect 150204 79872 150208 79928
rect 150208 79872 150264 79928
rect 150264 79872 150268 79928
rect 150204 79868 150268 79872
rect 150388 79928 150452 79932
rect 150388 79872 150392 79928
rect 150392 79872 150448 79928
rect 150448 79872 150452 79928
rect 150388 79868 150452 79872
rect 150940 79868 151004 79932
rect 151492 79868 151556 79932
rect 155724 80004 155788 80068
rect 159588 80140 159652 80204
rect 156276 80004 156340 80068
rect 149652 79732 149716 79796
rect 152228 79868 152292 79932
rect 153884 79928 153948 79932
rect 153884 79872 153888 79928
rect 153888 79872 153944 79928
rect 153944 79872 153948 79928
rect 153884 79868 153948 79872
rect 155356 79868 155420 79932
rect 156460 79868 156524 79932
rect 157196 79928 157260 79932
rect 157196 79872 157200 79928
rect 157200 79872 157256 79928
rect 157256 79872 157260 79928
rect 157196 79868 157260 79872
rect 157932 79868 157996 79932
rect 158300 79868 158364 79932
rect 152228 79792 152292 79796
rect 152228 79736 152232 79792
rect 152232 79736 152288 79792
rect 152288 79736 152292 79792
rect 152228 79732 152292 79736
rect 149836 79596 149900 79660
rect 151308 79656 151372 79660
rect 151308 79600 151322 79656
rect 151322 79600 151372 79656
rect 151308 79596 151372 79600
rect 153516 79732 153580 79796
rect 155356 79732 155420 79796
rect 157012 79732 157076 79796
rect 158852 79868 158916 79932
rect 160324 79928 160388 79932
rect 160324 79872 160328 79928
rect 160328 79872 160384 79928
rect 160384 79872 160388 79928
rect 160324 79868 160388 79872
rect 159036 79732 159100 79796
rect 154068 79596 154132 79660
rect 154252 79656 154316 79660
rect 154252 79600 154266 79656
rect 154266 79600 154316 79656
rect 154252 79596 154316 79600
rect 152596 79460 152660 79524
rect 153700 79460 153764 79524
rect 155724 79520 155788 79524
rect 155724 79464 155774 79520
rect 155774 79464 155788 79520
rect 155724 79460 155788 79464
rect 131988 79324 132052 79388
rect 152780 79324 152844 79388
rect 153884 79324 153948 79388
rect 167316 80140 167380 80204
rect 170628 80276 170692 80340
rect 161980 80004 162044 80068
rect 161428 79928 161492 79932
rect 161428 79872 161432 79928
rect 161432 79872 161488 79928
rect 161488 79872 161492 79928
rect 161428 79868 161492 79872
rect 160692 79792 160756 79796
rect 160692 79736 160742 79792
rect 160742 79736 160756 79792
rect 160692 79732 160756 79736
rect 156828 79596 156892 79660
rect 157748 79656 157812 79660
rect 157748 79600 157798 79656
rect 157798 79600 157812 79656
rect 157748 79596 157812 79600
rect 158116 79656 158180 79660
rect 158116 79600 158130 79656
rect 158130 79600 158180 79656
rect 158116 79596 158180 79600
rect 158668 79596 158732 79660
rect 157564 79460 157628 79524
rect 156828 79324 156892 79388
rect 125364 79188 125428 79252
rect 145236 79188 145300 79252
rect 148732 79188 148796 79252
rect 126652 79052 126716 79116
rect 138060 79052 138124 79116
rect 125180 78916 125244 78980
rect 145420 79052 145484 79116
rect 146708 79052 146772 79116
rect 147076 79052 147140 79116
rect 148180 79052 148244 79116
rect 149836 79052 149900 79116
rect 150020 79052 150084 79116
rect 160876 79656 160940 79660
rect 162164 79868 162228 79932
rect 163452 79868 163516 79932
rect 165476 80004 165540 80068
rect 165292 79928 165356 79932
rect 165292 79872 165296 79928
rect 165296 79872 165352 79928
rect 165352 79872 165356 79928
rect 165292 79868 165356 79872
rect 166396 80004 166460 80068
rect 164740 79792 164804 79796
rect 164740 79736 164754 79792
rect 164754 79736 164804 79792
rect 164740 79732 164804 79736
rect 165108 79732 165172 79796
rect 160876 79600 160926 79656
rect 160926 79600 160940 79656
rect 160876 79596 160940 79600
rect 162164 79596 162228 79660
rect 163084 79596 163148 79660
rect 163636 79596 163700 79660
rect 164188 79656 164252 79660
rect 164188 79600 164238 79656
rect 164238 79600 164252 79656
rect 164188 79596 164252 79600
rect 161612 79460 161676 79524
rect 162348 79460 162412 79524
rect 163268 79460 163332 79524
rect 164556 79460 164620 79524
rect 166580 79928 166644 79932
rect 166580 79872 166584 79928
rect 166584 79872 166640 79928
rect 166640 79872 166644 79928
rect 166580 79868 166644 79872
rect 166948 79928 167012 79932
rect 166948 79872 166952 79928
rect 166952 79872 167008 79928
rect 167008 79872 167012 79928
rect 166948 79868 167012 79872
rect 166028 79732 166092 79796
rect 167500 79732 167564 79796
rect 165844 79596 165908 79660
rect 168052 79928 168116 79932
rect 168052 79872 168056 79928
rect 168056 79872 168112 79928
rect 168112 79872 168116 79928
rect 168052 79868 168116 79872
rect 168236 79906 168240 79932
rect 168240 79906 168296 79932
rect 168296 79906 168300 79932
rect 168236 79868 168300 79906
rect 168604 80004 168668 80068
rect 170260 80140 170324 80204
rect 172836 80140 172900 80204
rect 169340 79732 169404 79796
rect 170996 79868 171060 79932
rect 171548 79928 171612 79932
rect 171548 79872 171552 79928
rect 171552 79872 171608 79928
rect 171608 79872 171612 79928
rect 171548 79868 171612 79872
rect 171732 79868 171796 79932
rect 169708 79732 169772 79796
rect 169892 79732 169956 79796
rect 171180 79732 171244 79796
rect 172100 79732 172164 79796
rect 167868 79596 167932 79660
rect 166764 79460 166828 79524
rect 167316 79460 167380 79524
rect 167684 79460 167748 79524
rect 169156 79596 169220 79660
rect 170076 79596 170140 79660
rect 171364 79596 171428 79660
rect 169524 79460 169588 79524
rect 170628 79460 170692 79524
rect 159956 79324 160020 79388
rect 170444 79324 170508 79388
rect 164004 79188 164068 79252
rect 164924 79188 164988 79252
rect 166212 79188 166276 79252
rect 173020 79868 173084 79932
rect 175596 80140 175660 80204
rect 176332 80140 176396 80204
rect 173020 79732 173084 79796
rect 173572 79732 173636 79796
rect 174860 79868 174924 79932
rect 175044 79868 175108 79932
rect 175596 79868 175660 79932
rect 176148 79868 176212 79932
rect 176332 79928 176396 79932
rect 176332 79872 176336 79928
rect 176336 79872 176392 79928
rect 176392 79872 176396 79928
rect 176332 79868 176396 79872
rect 174124 79732 174188 79796
rect 174676 79732 174740 79796
rect 175964 79732 176028 79796
rect 186268 80004 186332 80068
rect 177068 79868 177132 79932
rect 177620 79868 177684 79932
rect 176884 79732 176948 79796
rect 173388 79596 173452 79660
rect 174308 79596 174372 79660
rect 175780 79596 175844 79660
rect 172652 79460 172716 79524
rect 175412 79460 175476 79524
rect 177068 79460 177132 79524
rect 177804 79460 177868 79524
rect 180932 79460 180996 79524
rect 171916 79188 171980 79252
rect 175228 79188 175292 79252
rect 175964 79188 176028 79252
rect 193996 79324 194060 79388
rect 190868 79188 190932 79252
rect 160692 79052 160756 79116
rect 162532 79052 162596 79116
rect 166948 79052 167012 79116
rect 167868 79052 167932 79116
rect 168972 79052 169036 79116
rect 170812 79052 170876 79116
rect 140452 78916 140516 78980
rect 142108 78916 142172 78980
rect 142660 78916 142724 78980
rect 143212 78916 143276 78980
rect 145604 78916 145668 78980
rect 170996 78916 171060 78980
rect 173204 79052 173268 79116
rect 172100 78916 172164 78980
rect 176516 78916 176580 78980
rect 179460 78976 179524 78980
rect 179460 78920 179510 78976
rect 179510 78920 179524 78976
rect 179460 78916 179524 78920
rect 180748 78916 180812 78980
rect 198964 78916 199028 78980
rect 199332 78916 199396 78980
rect 124076 78780 124140 78844
rect 130884 78644 130948 78708
rect 124812 78508 124876 78572
rect 132908 78568 132972 78572
rect 132908 78512 132922 78568
rect 132922 78512 132972 78568
rect 132908 78508 132972 78512
rect 133460 78508 133524 78572
rect 135852 78508 135916 78572
rect 137140 78508 137204 78572
rect 138060 78568 138124 78572
rect 138060 78512 138110 78568
rect 138110 78512 138124 78568
rect 138060 78508 138124 78512
rect 139348 78644 139412 78708
rect 143396 78644 143460 78708
rect 148916 78780 148980 78844
rect 151492 78644 151556 78708
rect 158116 78704 158180 78708
rect 158116 78648 158166 78704
rect 158166 78648 158180 78704
rect 158116 78644 158180 78648
rect 158484 78704 158548 78708
rect 158484 78648 158534 78704
rect 158534 78648 158548 78704
rect 158484 78644 158548 78648
rect 159588 78644 159652 78708
rect 168236 78704 168300 78708
rect 168236 78648 168286 78704
rect 168286 78648 168300 78704
rect 168236 78644 168300 78648
rect 152412 78568 152476 78572
rect 152412 78512 152426 78568
rect 152426 78512 152476 78568
rect 128124 78372 128188 78436
rect 152412 78508 152476 78512
rect 154068 78568 154132 78572
rect 154068 78512 154082 78568
rect 154082 78512 154132 78568
rect 154068 78508 154132 78512
rect 154436 78568 154500 78572
rect 154436 78512 154486 78568
rect 154486 78512 154500 78568
rect 154436 78508 154500 78512
rect 155724 78508 155788 78572
rect 171916 78508 171980 78572
rect 173388 78508 173452 78572
rect 174860 78568 174924 78572
rect 174860 78512 174874 78568
rect 174874 78512 174924 78568
rect 174860 78508 174924 78512
rect 177620 78508 177684 78572
rect 126836 78236 126900 78300
rect 135484 78236 135548 78300
rect 142476 78372 142540 78436
rect 150756 78372 150820 78436
rect 156644 78372 156708 78436
rect 159036 78372 159100 78436
rect 173020 78372 173084 78436
rect 187924 78372 187988 78436
rect 148364 78236 148428 78300
rect 149100 78236 149164 78300
rect 152412 78236 152476 78300
rect 168604 78236 168668 78300
rect 171548 78236 171612 78300
rect 131804 77964 131868 78028
rect 151124 78100 151188 78164
rect 152964 78100 153028 78164
rect 156276 78160 156340 78164
rect 156276 78104 156326 78160
rect 156326 78104 156340 78160
rect 156276 78100 156340 78104
rect 175964 78160 176028 78164
rect 175964 78104 176014 78160
rect 176014 78104 176028 78160
rect 175964 78100 176028 78104
rect 176332 78236 176396 78300
rect 198964 78100 199028 78164
rect 147444 77964 147508 78028
rect 166396 77964 166460 78028
rect 136036 77828 136100 77892
rect 152780 77828 152844 77892
rect 153700 77828 153764 77892
rect 155540 77828 155604 77892
rect 157012 77828 157076 77892
rect 158300 77828 158364 77892
rect 177068 77828 177132 77892
rect 138612 77692 138676 77756
rect 140636 77692 140700 77756
rect 148548 77692 148612 77756
rect 149468 77692 149532 77756
rect 126468 77556 126532 77620
rect 130332 77420 130396 77484
rect 138244 77556 138308 77620
rect 156460 77556 156524 77620
rect 165108 77616 165172 77620
rect 165108 77560 165122 77616
rect 165122 77560 165172 77616
rect 165108 77556 165172 77560
rect 170996 77556 171060 77620
rect 171732 77556 171796 77620
rect 139164 77420 139228 77484
rect 140820 77480 140884 77484
rect 140820 77424 140870 77480
rect 140870 77424 140884 77480
rect 140820 77420 140884 77424
rect 174492 77556 174556 77620
rect 134748 77284 134812 77348
rect 140268 77284 140332 77348
rect 140820 77284 140884 77348
rect 160876 77344 160940 77348
rect 160876 77288 160890 77344
rect 160890 77288 160940 77344
rect 134932 77148 134996 77212
rect 160876 77284 160940 77288
rect 161060 77344 161124 77348
rect 187924 77828 187988 77892
rect 161060 77288 161110 77344
rect 161110 77288 161124 77344
rect 161060 77284 161124 77288
rect 143028 77148 143092 77212
rect 176148 77148 176212 77212
rect 178908 77148 178972 77212
rect 180012 77208 180076 77212
rect 180012 77152 180062 77208
rect 180062 77152 180076 77208
rect 180012 77148 180076 77152
rect 146892 77012 146956 77076
rect 191972 77012 192036 77076
rect 169340 76876 169404 76940
rect 174860 76876 174924 76940
rect 148180 76740 148244 76804
rect 178540 76740 178604 76804
rect 134380 76604 134444 76668
rect 153884 76664 153948 76668
rect 153884 76608 153934 76664
rect 153934 76608 153948 76664
rect 153884 76604 153948 76608
rect 170260 76604 170324 76668
rect 191604 76604 191668 76668
rect 162532 76468 162596 76532
rect 170812 76468 170876 76532
rect 183692 76332 183756 76396
rect 163268 76120 163332 76124
rect 163268 76064 163318 76120
rect 163318 76064 163332 76120
rect 163268 76060 163332 76064
rect 165476 76060 165540 76124
rect 134012 75924 134076 75988
rect 135668 75924 135732 75988
rect 135852 75984 135916 75988
rect 135852 75928 135902 75984
rect 135902 75928 135916 75984
rect 135852 75924 135916 75928
rect 148732 75924 148796 75988
rect 162716 75924 162780 75988
rect 163452 75924 163516 75988
rect 166396 75984 166460 75988
rect 166396 75928 166446 75984
rect 166446 75928 166460 75984
rect 166396 75924 166460 75928
rect 166580 75924 166644 75988
rect 167684 75924 167748 75988
rect 173572 75924 173636 75988
rect 135484 75788 135548 75852
rect 139348 75652 139412 75716
rect 152964 75652 153028 75716
rect 141004 75516 141068 75580
rect 174676 75576 174740 75580
rect 174676 75520 174726 75576
rect 174726 75520 174740 75576
rect 174676 75516 174740 75520
rect 175596 75516 175660 75580
rect 193260 75516 193324 75580
rect 145604 75380 145668 75444
rect 196388 75380 196452 75444
rect 171180 75244 171244 75308
rect 170996 75108 171060 75172
rect 148364 74972 148428 75036
rect 181116 74972 181180 75036
rect 189028 74972 189092 75036
rect 137508 74836 137572 74900
rect 144684 74700 144748 74764
rect 122788 74564 122852 74628
rect 118556 74428 118620 74492
rect 156460 74428 156524 74492
rect 122788 74292 122852 74356
rect 193812 74292 193876 74356
rect 134380 74156 134444 74220
rect 183508 74156 183572 74220
rect 139716 74020 139780 74084
rect 177068 74020 177132 74084
rect 187740 74020 187804 74084
rect 140820 73884 140884 73948
rect 145052 73884 145116 73948
rect 192524 73884 192588 73948
rect 122604 73748 122668 73812
rect 181300 73748 181364 73812
rect 158484 73612 158548 73676
rect 179828 73612 179892 73676
rect 122420 73068 122484 73132
rect 156828 73068 156892 73132
rect 139532 72932 139596 72996
rect 183140 72932 183204 72996
rect 151124 72796 151188 72860
rect 196572 72796 196636 72860
rect 149100 72660 149164 72724
rect 149468 72660 149532 72724
rect 150020 72524 150084 72588
rect 145420 72252 145484 72316
rect 184980 71708 185044 71772
rect 118188 71572 118252 71636
rect 152412 71572 152476 71636
rect 173572 71572 173636 71636
rect 197492 71572 197556 71636
rect 149652 71436 149716 71500
rect 184060 71436 184124 71500
rect 145052 71300 145116 71364
rect 187740 71164 187804 71228
rect 144132 71028 144196 71092
rect 197492 71028 197556 71092
rect 198044 71028 198108 71092
rect 142108 70408 142172 70412
rect 142108 70352 142122 70408
rect 142122 70352 142172 70408
rect 142108 70348 142172 70352
rect 122236 70212 122300 70276
rect 175964 70212 176028 70276
rect 201356 70212 201420 70276
rect 148732 70076 148796 70140
rect 182772 70076 182836 70140
rect 144500 69940 144564 70004
rect 178356 69940 178420 70004
rect 201356 69532 201420 69596
rect 144684 68852 144748 68916
rect 145604 68852 145668 68916
rect 182956 68912 183020 68916
rect 182956 68856 183006 68912
rect 183006 68856 183020 68912
rect 182956 68852 183020 68856
rect 198780 68852 198844 68916
rect 176148 68716 176212 68780
rect 144316 68580 144380 68644
rect 148548 68308 148612 68372
rect 135668 67492 135732 67556
rect 189028 67492 189092 67556
rect 155540 67356 155604 67420
rect 151492 67220 151556 67284
rect 178172 67220 178236 67284
rect 148180 67084 148244 67148
rect 133644 66812 133708 66876
rect 146892 66812 146956 66876
rect 162164 66676 162228 66740
rect 137508 66132 137572 66196
rect 153884 66132 153948 66196
rect 160692 65996 160756 66060
rect 171916 65724 171980 65788
rect 189396 65724 189460 65788
rect 173756 65452 173820 65516
rect 195100 65452 195164 65516
rect 142108 64968 142172 64972
rect 142108 64912 142122 64968
rect 142122 64912 142172 64968
rect 142108 64908 142172 64912
rect 174676 64772 174740 64836
rect 197860 64772 197924 64836
rect 142108 64636 142172 64700
rect 172100 64636 172164 64700
rect 187004 64636 187068 64700
rect 187004 64228 187068 64292
rect 197860 64092 197924 64156
rect 138612 63412 138676 63476
rect 166212 63412 166276 63476
rect 149468 63276 149532 63340
rect 154068 63140 154132 63204
rect 155724 63004 155788 63068
rect 174860 62868 174924 62932
rect 197308 62868 197372 62932
rect 187188 62052 187252 62116
rect 196020 62112 196084 62116
rect 196020 62056 196070 62112
rect 196070 62056 196084 62112
rect 196020 62052 196084 62056
rect 157012 61916 157076 61980
rect 164924 61780 164988 61844
rect 149836 61644 149900 61708
rect 165108 60556 165172 60620
rect 176332 60420 176396 60484
rect 200988 59876 201052 59940
rect 188292 59332 188356 59396
rect 167500 59196 167564 59260
rect 154252 59060 154316 59124
rect 157932 58788 157996 58852
rect 162348 58652 162412 58716
rect 120764 57972 120828 58036
rect 134380 57836 134444 57900
rect 152780 57836 152844 57900
rect 138428 57700 138492 57764
rect 156644 57564 156708 57628
rect 160876 57428 160940 57492
rect 165292 57292 165356 57356
rect 175044 57156 175108 57220
rect 200804 57156 200868 57220
rect 167684 56476 167748 56540
rect 158852 56340 158916 56404
rect 163268 56204 163332 56268
rect 176516 56068 176580 56132
rect 200620 56068 200684 56132
rect 201356 56068 201420 56132
rect 172284 55932 172348 55996
rect 201356 55796 201420 55860
rect 142108 55312 142172 55316
rect 142108 55256 142122 55312
rect 142122 55256 142172 55312
rect 142108 55252 142172 55256
rect 138244 55116 138308 55180
rect 163452 55116 163516 55180
rect 201724 55176 201788 55180
rect 201724 55120 201738 55176
rect 201738 55120 201788 55176
rect 201724 55116 201788 55120
rect 142108 54980 142172 55044
rect 158116 54980 158180 55044
rect 161060 54844 161124 54908
rect 166396 53756 166460 53820
rect 162532 53620 162596 53684
rect 154436 53484 154500 53548
rect 182588 53348 182652 53412
rect 134196 52396 134260 52460
rect 167868 52396 167932 52460
rect 163636 52260 163700 52324
rect 134012 50900 134076 50964
rect 165476 50900 165540 50964
rect 203012 50960 203076 50964
rect 203012 50904 203062 50960
rect 203062 50904 203076 50960
rect 203012 50900 203076 50904
rect 158300 50764 158364 50828
rect 144684 50628 144748 50692
rect 135484 49540 135548 49604
rect 166580 49540 166644 49604
rect 162716 49404 162780 49468
rect 159036 49268 159100 49332
rect 190500 48996 190564 49060
rect 135852 48180 135916 48244
rect 169340 48180 169404 48244
rect 161244 48044 161308 48108
rect 137692 46820 137756 46884
rect 168052 46820 168116 46884
rect 201540 46140 201604 46204
rect 142108 45656 142172 45660
rect 142108 45600 142122 45656
rect 142122 45600 142172 45656
rect 142108 45596 142172 45600
rect 192340 45596 192404 45660
rect 142108 45520 142172 45524
rect 142108 45464 142122 45520
rect 142122 45464 142172 45520
rect 142108 45460 142172 45464
rect 146708 44916 146772 44980
rect 151124 44780 151188 44844
rect 138060 44100 138124 44164
rect 166764 44100 166828 44164
rect 169524 43964 169588 44028
rect 149284 42060 149348 42124
rect 152964 40564 153028 40628
rect 133460 36484 133524 36548
rect 170996 36484 171060 36548
rect 142108 36076 142172 36140
rect 142292 35804 142356 35868
rect 134932 33764 134996 33828
rect 148916 32404 148980 32468
rect 120580 31724 120644 31788
rect 145420 26964 145484 27028
rect 152412 26828 152476 26892
rect 142108 26344 142172 26348
rect 142108 26288 142122 26344
rect 142122 26288 142172 26344
rect 142108 26284 142172 26288
rect 142108 26208 142172 26212
rect 142108 26152 142122 26208
rect 142122 26152 142172 26208
rect 142108 26148 142172 26152
rect 144500 21252 144564 21316
rect 116532 19348 116596 19412
rect 149652 18532 149716 18596
rect 142292 16628 142356 16692
rect 142108 16356 142172 16420
rect 144316 15812 144380 15876
rect 158484 11596 158548 11660
rect 142108 7032 142172 7036
rect 142108 6976 142122 7032
rect 142122 6976 142172 7032
rect 142108 6972 142172 6976
rect 142108 6896 142172 6900
rect 142108 6840 142122 6896
rect 142122 6840 142172 6896
rect 142108 6836 142172 6840
rect 144132 4796 144196 4860
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 111563 265164 111629 265165
rect 111563 265100 111564 265164
rect 111628 265100 111629 265164
rect 111563 265099 111629 265100
rect 111379 261084 111445 261085
rect 111379 261020 111380 261084
rect 111444 261020 111445 261084
rect 111379 261019 111445 261020
rect 111195 260948 111261 260949
rect 111195 260884 111196 260948
rect 111260 260884 111261 260948
rect 111195 260883 111261 260884
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 111198 146029 111258 260883
rect 111195 146028 111261 146029
rect 111195 145964 111196 146028
rect 111260 145964 111261 146028
rect 111195 145963 111261 145964
rect 111382 143309 111442 261019
rect 111566 146165 111626 265099
rect 113035 265028 113101 265029
rect 113035 264964 113036 265028
rect 113100 264964 113101 265028
rect 113035 264963 113101 264964
rect 112851 263668 112917 263669
rect 112851 263604 112852 263668
rect 112916 263604 112917 263668
rect 112851 263603 112917 263604
rect 112667 262716 112733 262717
rect 112667 262652 112668 262716
rect 112732 262652 112733 262716
rect 112667 262651 112733 262652
rect 111563 146164 111629 146165
rect 111563 146100 111564 146164
rect 111628 146100 111629 146164
rect 111563 146099 111629 146100
rect 112670 144533 112730 262651
rect 112667 144532 112733 144533
rect 112667 144468 112668 144532
rect 112732 144468 112733 144532
rect 112667 144467 112733 144468
rect 112854 144397 112914 263603
rect 112851 144396 112917 144397
rect 112851 144332 112852 144396
rect 112916 144332 112917 144396
rect 112851 144331 112917 144332
rect 113038 143853 113098 264963
rect 114139 262988 114205 262989
rect 114139 262924 114140 262988
rect 114204 262924 114205 262988
rect 114139 262923 114205 262924
rect 113955 262580 114021 262581
rect 113955 262516 113956 262580
rect 114020 262516 114021 262580
rect 113955 262515 114021 262516
rect 113771 259724 113837 259725
rect 113771 259660 113772 259724
rect 113836 259660 113837 259724
rect 113771 259659 113837 259660
rect 113774 145893 113834 259659
rect 113771 145892 113837 145893
rect 113771 145828 113772 145892
rect 113836 145828 113837 145892
rect 113771 145827 113837 145828
rect 113958 145621 114018 262515
rect 114142 145757 114202 262923
rect 114294 259954 114914 295398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 115611 262852 115677 262853
rect 115611 262788 115612 262852
rect 115676 262788 115677 262852
rect 115611 262787 115677 262788
rect 115427 262308 115493 262309
rect 115427 262244 115428 262308
rect 115492 262244 115493 262308
rect 115427 262243 115493 262244
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114139 145756 114205 145757
rect 114139 145692 114140 145756
rect 114204 145692 114205 145756
rect 114139 145691 114205 145692
rect 113955 145620 114021 145621
rect 113955 145556 113956 145620
rect 114020 145556 114021 145620
rect 113955 145555 114021 145556
rect 113035 143852 113101 143853
rect 113035 143788 113036 143852
rect 113100 143788 113101 143852
rect 113035 143787 113101 143788
rect 111379 143308 111445 143309
rect 111379 143244 111380 143308
rect 111444 143244 111445 143308
rect 111379 143243 111445 143244
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 115954 114914 151398
rect 115430 146301 115490 262243
rect 115427 146300 115493 146301
rect 115427 146236 115428 146300
rect 115492 146236 115493 146300
rect 115427 146235 115493 146236
rect 115614 143989 115674 262787
rect 116715 262444 116781 262445
rect 116715 262380 116716 262444
rect 116780 262380 116781 262444
rect 116715 262379 116781 262380
rect 115795 259588 115861 259589
rect 115795 259524 115796 259588
rect 115860 259524 115861 259588
rect 115795 259523 115861 259524
rect 115611 143988 115677 143989
rect 115611 143924 115612 143988
rect 115676 143924 115677 143988
rect 115611 143923 115677 143924
rect 115798 141405 115858 259523
rect 116718 144125 116778 262379
rect 118794 262000 119414 263898
rect 119843 263940 119909 263941
rect 119843 263876 119844 263940
rect 119908 263876 119909 263940
rect 119843 263875 119909 263876
rect 117083 260404 117149 260405
rect 117083 260340 117084 260404
rect 117148 260340 117149 260404
rect 117083 260339 117149 260340
rect 116899 259996 116965 259997
rect 116899 259932 116900 259996
rect 116964 259932 116965 259996
rect 116899 259931 116965 259932
rect 116715 144124 116781 144125
rect 116715 144060 116716 144124
rect 116780 144060 116781 144124
rect 116715 144059 116781 144060
rect 116902 141541 116962 259931
rect 117086 141813 117146 260339
rect 118371 260132 118437 260133
rect 118371 260068 118372 260132
rect 118436 260068 118437 260132
rect 118371 260067 118437 260068
rect 118187 259860 118253 259861
rect 118187 259796 118188 259860
rect 118252 259796 118253 259860
rect 118187 259795 118253 259796
rect 118190 144805 118250 259795
rect 118187 144804 118253 144805
rect 118187 144740 118188 144804
rect 118252 144740 118253 144804
rect 118187 144739 118253 144740
rect 118187 144260 118253 144261
rect 118187 144196 118188 144260
rect 118252 144196 118253 144260
rect 118187 144195 118253 144196
rect 117083 141812 117149 141813
rect 117083 141748 117084 141812
rect 117148 141748 117149 141812
rect 117083 141747 117149 141748
rect 116899 141540 116965 141541
rect 116899 141476 116900 141540
rect 116964 141476 116965 141540
rect 116899 141475 116965 141476
rect 115795 141404 115861 141405
rect 115795 141340 115796 141404
rect 115860 141340 115861 141404
rect 115795 141339 115861 141340
rect 116531 140452 116597 140453
rect 116531 140388 116532 140452
rect 116596 140388 116597 140452
rect 116531 140387 116597 140388
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 116534 19413 116594 140387
rect 118190 71637 118250 144195
rect 118374 141677 118434 260067
rect 118555 196620 118621 196621
rect 118555 196556 118556 196620
rect 118620 196556 118621 196620
rect 118555 196555 118621 196556
rect 118371 141676 118437 141677
rect 118371 141612 118372 141676
rect 118436 141612 118437 141676
rect 118371 141611 118437 141612
rect 118558 74493 118618 196555
rect 118794 192454 119414 198000
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 119846 142901 119906 263875
rect 121315 263804 121381 263805
rect 121315 263740 121316 263804
rect 121380 263740 121381 263804
rect 121315 263739 121381 263740
rect 121131 260268 121197 260269
rect 121131 260204 121132 260268
rect 121196 260204 121197 260268
rect 121131 260203 121197 260204
rect 120763 144940 120829 144941
rect 120763 144876 120764 144940
rect 120828 144876 120829 144940
rect 120763 144875 120829 144876
rect 119843 142900 119909 142901
rect 119843 142836 119844 142900
rect 119908 142836 119909 142900
rect 119843 142835 119909 142836
rect 120579 140588 120645 140589
rect 120579 140524 120580 140588
rect 120644 140524 120645 140588
rect 120579 140523 120645 140524
rect 119291 139908 119357 139909
rect 119291 139844 119292 139908
rect 119356 139844 119357 139908
rect 119291 139843 119357 139844
rect 119294 84285 119354 139843
rect 119291 84284 119357 84285
rect 119291 84220 119292 84284
rect 119356 84220 119357 84284
rect 119291 84219 119357 84220
rect 118555 74492 118621 74493
rect 118555 74428 118556 74492
rect 118620 74428 118621 74492
rect 118555 74427 118621 74428
rect 118187 71636 118253 71637
rect 118187 71572 118188 71636
rect 118252 71572 118253 71636
rect 118187 71571 118253 71572
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 116531 19412 116597 19413
rect 116531 19348 116532 19412
rect 116596 19348 116597 19412
rect 116531 19347 116597 19348
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 12454 119414 47898
rect 120582 31789 120642 140523
rect 120766 58037 120826 144875
rect 121134 143173 121194 260203
rect 121131 143172 121197 143173
rect 121131 143108 121132 143172
rect 121196 143108 121197 143172
rect 121131 143107 121197 143108
rect 121318 143037 121378 263739
rect 123294 262000 123914 268398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 262000 128414 272898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 262000 132914 277398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 262000 137414 281898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 262000 141914 286398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 262000 146414 290898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 262000 150914 295398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 262000 155414 263898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 262000 159914 268398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 262000 164414 272898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 262000 168914 277398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 262000 173414 281898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 262000 177914 286398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 262000 182414 290898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 262000 186914 295398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 189027 278084 189093 278085
rect 189027 278020 189028 278084
rect 189092 278020 189093 278084
rect 189027 278019 189093 278020
rect 189030 277541 189090 278019
rect 189027 277540 189093 277541
rect 189027 277476 189028 277540
rect 189092 277476 189093 277540
rect 189027 277475 189093 277476
rect 186083 259588 186149 259589
rect 186083 259524 186084 259588
rect 186148 259524 186149 259588
rect 186083 259523 186149 259524
rect 124208 255454 124528 255486
rect 124208 255218 124250 255454
rect 124486 255218 124528 255454
rect 124208 255134 124528 255218
rect 124208 254898 124250 255134
rect 124486 254898 124528 255134
rect 124208 254866 124528 254898
rect 154928 255454 155248 255486
rect 154928 255218 154970 255454
rect 155206 255218 155248 255454
rect 154928 255134 155248 255218
rect 154928 254898 154970 255134
rect 155206 254898 155248 255134
rect 154928 254866 155248 254898
rect 185648 255454 185968 255486
rect 185648 255218 185690 255454
rect 185926 255218 185968 255454
rect 185648 255134 185968 255218
rect 185648 254898 185690 255134
rect 185926 254898 185968 255134
rect 185648 254866 185968 254898
rect 139568 223954 139888 223986
rect 139568 223718 139610 223954
rect 139846 223718 139888 223954
rect 139568 223634 139888 223718
rect 139568 223398 139610 223634
rect 139846 223398 139888 223634
rect 139568 223366 139888 223398
rect 170288 223954 170608 223986
rect 170288 223718 170330 223954
rect 170566 223718 170608 223954
rect 170288 223634 170608 223718
rect 170288 223398 170330 223634
rect 170566 223398 170608 223634
rect 170288 223366 170608 223398
rect 124208 219454 124528 219486
rect 124208 219218 124250 219454
rect 124486 219218 124528 219454
rect 124208 219134 124528 219218
rect 124208 218898 124250 219134
rect 124486 218898 124528 219134
rect 124208 218866 124528 218898
rect 154928 219454 155248 219486
rect 154928 219218 154970 219454
rect 155206 219218 155248 219454
rect 154928 219134 155248 219218
rect 154928 218898 154970 219134
rect 155206 218898 155248 219134
rect 154928 218866 155248 218898
rect 185648 219454 185968 219486
rect 185648 219218 185690 219454
rect 185926 219218 185968 219454
rect 185648 219134 185968 219218
rect 185648 218898 185690 219134
rect 185926 218898 185968 219134
rect 185648 218866 185968 218898
rect 186086 212533 186146 259523
rect 186083 212532 186149 212533
rect 186083 212468 186084 212532
rect 186148 212468 186149 212532
rect 186083 212467 186149 212468
rect 187187 212532 187253 212533
rect 187187 212468 187188 212532
rect 187252 212468 187253 212532
rect 187187 212467 187253 212468
rect 141555 200700 141621 200701
rect 141555 200636 141556 200700
rect 141620 200636 141621 200700
rect 141555 200635 141621 200636
rect 136587 200564 136653 200565
rect 136587 200500 136588 200564
rect 136652 200500 136653 200564
rect 136587 200499 136653 200500
rect 133643 200156 133709 200157
rect 133643 200092 133644 200156
rect 133708 200092 133709 200156
rect 133643 200091 133709 200092
rect 133646 199885 133706 200091
rect 133091 199884 133157 199885
rect 133091 199820 133092 199884
rect 133156 199820 133157 199884
rect 133091 199819 133157 199820
rect 133643 199884 133709 199885
rect 133643 199820 133644 199884
rect 133708 199820 133709 199884
rect 133643 199819 133709 199820
rect 134747 199884 134813 199885
rect 134747 199820 134748 199884
rect 134812 199820 134813 199884
rect 134747 199819 134813 199820
rect 136035 199884 136101 199885
rect 136035 199820 136036 199884
rect 136100 199820 136101 199884
rect 136035 199819 136101 199820
rect 122603 199476 122669 199477
rect 122603 199412 122604 199476
rect 122668 199412 122669 199476
rect 122603 199411 122669 199412
rect 122419 147796 122485 147797
rect 122419 147732 122420 147796
rect 122484 147732 122485 147796
rect 122419 147731 122485 147732
rect 121315 143036 121381 143037
rect 121315 142972 121316 143036
rect 121380 142972 121381 143036
rect 121315 142971 121381 142972
rect 122235 140180 122301 140181
rect 122235 140116 122236 140180
rect 122300 140116 122301 140180
rect 122235 140115 122301 140116
rect 122051 139364 122117 139365
rect 122051 139300 122052 139364
rect 122116 139300 122117 139364
rect 122051 139299 122117 139300
rect 122054 128370 122114 139299
rect 122238 138005 122298 140115
rect 122235 138004 122301 138005
rect 122235 137940 122236 138004
rect 122300 137940 122301 138004
rect 122235 137939 122301 137940
rect 122054 128310 122298 128370
rect 122238 70277 122298 128310
rect 122422 73133 122482 147731
rect 122606 73813 122666 199411
rect 133094 198750 133154 199819
rect 133094 198690 133338 198750
rect 130883 198524 130949 198525
rect 130883 198460 130884 198524
rect 130948 198460 130949 198524
rect 130883 198459 130949 198460
rect 125363 198388 125429 198389
rect 125363 198324 125364 198388
rect 125428 198324 125429 198388
rect 125363 198323 125429 198324
rect 125179 198252 125245 198253
rect 125179 198188 125180 198252
rect 125244 198188 125245 198252
rect 125179 198187 125245 198188
rect 124995 198116 125061 198117
rect 124995 198052 124996 198116
rect 125060 198052 125061 198116
rect 124995 198051 125061 198052
rect 123294 196954 123914 198000
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 124075 195260 124141 195261
rect 124075 195196 124076 195260
rect 124140 195196 124141 195260
rect 124075 195195 124141 195196
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 122971 142220 123037 142221
rect 122971 142156 122972 142220
rect 123036 142156 123037 142220
rect 122971 142155 123037 142156
rect 122787 138004 122853 138005
rect 122787 137940 122788 138004
rect 122852 137940 122853 138004
rect 122787 137939 122853 137940
rect 122790 128485 122850 137939
rect 122787 128484 122853 128485
rect 122787 128420 122788 128484
rect 122852 128420 122853 128484
rect 122787 128419 122853 128420
rect 122787 123180 122853 123181
rect 122787 123116 122788 123180
rect 122852 123116 122853 123180
rect 122787 123115 122853 123116
rect 122790 122501 122850 123115
rect 122787 122500 122853 122501
rect 122787 122436 122788 122500
rect 122852 122436 122853 122500
rect 122787 122435 122853 122436
rect 122787 113524 122853 113525
rect 122787 113460 122788 113524
rect 122852 113460 122853 113524
rect 122787 113459 122853 113460
rect 122790 112845 122850 113459
rect 122787 112844 122853 112845
rect 122787 112780 122788 112844
rect 122852 112780 122853 112844
rect 122787 112779 122853 112780
rect 122787 103868 122853 103869
rect 122787 103804 122788 103868
rect 122852 103804 122853 103868
rect 122787 103803 122853 103804
rect 122790 103189 122850 103803
rect 122787 103188 122853 103189
rect 122787 103124 122788 103188
rect 122852 103124 122853 103188
rect 122787 103123 122853 103124
rect 122787 94212 122853 94213
rect 122787 94148 122788 94212
rect 122852 94148 122853 94212
rect 122787 94147 122853 94148
rect 122790 93533 122850 94147
rect 122787 93532 122853 93533
rect 122787 93468 122788 93532
rect 122852 93468 122853 93532
rect 122787 93467 122853 93468
rect 122787 89724 122853 89725
rect 122787 89660 122788 89724
rect 122852 89660 122853 89724
rect 122787 89659 122853 89660
rect 122790 80341 122850 89659
rect 122787 80340 122853 80341
rect 122787 80276 122788 80340
rect 122852 80276 122853 80340
rect 122787 80275 122853 80276
rect 122974 80069 123034 142155
rect 123294 142000 123914 160398
rect 122971 80068 123037 80069
rect 122971 80004 122972 80068
rect 123036 80004 123037 80068
rect 122971 80003 123037 80004
rect 124078 78845 124138 195195
rect 124811 194172 124877 194173
rect 124811 194108 124812 194172
rect 124876 194108 124877 194172
rect 124811 194107 124877 194108
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 124075 78844 124141 78845
rect 124075 78780 124076 78844
rect 124140 78780 124141 78844
rect 124075 78779 124141 78780
rect 124814 78573 124874 194107
rect 124998 80885 125058 198051
rect 124995 80884 125061 80885
rect 124995 80820 124996 80884
rect 125060 80820 125061 80884
rect 124995 80819 125061 80820
rect 125182 78981 125242 198187
rect 125366 79253 125426 198323
rect 130699 197572 130765 197573
rect 130699 197508 130700 197572
rect 130764 197508 130765 197572
rect 130699 197507 130765 197508
rect 126651 197436 126717 197437
rect 126651 197372 126652 197436
rect 126716 197372 126717 197436
rect 126651 197371 126717 197372
rect 130515 197436 130581 197437
rect 130515 197372 130516 197436
rect 130580 197372 130581 197436
rect 130515 197371 130581 197372
rect 126467 195532 126533 195533
rect 126467 195468 126468 195532
rect 126532 195468 126533 195532
rect 126467 195467 126533 195468
rect 126283 139364 126349 139365
rect 126283 139300 126284 139364
rect 126348 139300 126349 139364
rect 126283 139299 126349 139300
rect 126286 80341 126346 139299
rect 126283 80340 126349 80341
rect 126283 80276 126284 80340
rect 126348 80276 126349 80340
rect 126283 80275 126349 80276
rect 125363 79252 125429 79253
rect 125363 79188 125364 79252
rect 125428 79188 125429 79252
rect 125363 79187 125429 79188
rect 125179 78980 125245 78981
rect 125179 78916 125180 78980
rect 125244 78916 125245 78980
rect 125179 78915 125245 78916
rect 124811 78572 124877 78573
rect 124811 78508 124812 78572
rect 124876 78508 124877 78572
rect 124811 78507 124877 78508
rect 122787 74628 122853 74629
rect 122787 74564 122788 74628
rect 122852 74564 122853 74628
rect 122787 74563 122853 74564
rect 122790 74357 122850 74563
rect 122787 74356 122853 74357
rect 122787 74292 122788 74356
rect 122852 74292 122853 74356
rect 122787 74291 122853 74292
rect 122603 73812 122669 73813
rect 122603 73748 122604 73812
rect 122668 73748 122669 73812
rect 122603 73747 122669 73748
rect 122419 73132 122485 73133
rect 122419 73068 122420 73132
rect 122484 73068 122485 73132
rect 122419 73067 122485 73068
rect 122235 70276 122301 70277
rect 122235 70212 122236 70276
rect 122300 70212 122301 70276
rect 122235 70211 122301 70212
rect 120763 58036 120829 58037
rect 120763 57972 120764 58036
rect 120828 57972 120829 58036
rect 120763 57971 120829 57972
rect 123294 52954 123914 78000
rect 126470 77621 126530 195467
rect 126654 79117 126714 197371
rect 126835 197300 126901 197301
rect 126835 197236 126836 197300
rect 126900 197236 126901 197300
rect 126835 197235 126901 197236
rect 126651 79116 126717 79117
rect 126651 79052 126652 79116
rect 126716 79052 126717 79116
rect 126651 79051 126717 79052
rect 126838 78301 126898 197235
rect 128123 195804 128189 195805
rect 128123 195740 128124 195804
rect 128188 195740 128189 195804
rect 128123 195739 128189 195740
rect 127939 139364 128005 139365
rect 127939 139300 127940 139364
rect 128004 139300 128005 139364
rect 127939 139299 128005 139300
rect 127942 81021 128002 139299
rect 127939 81020 128005 81021
rect 127939 80956 127940 81020
rect 128004 80956 128005 81020
rect 127939 80955 128005 80956
rect 128126 78437 128186 195739
rect 130331 194036 130397 194037
rect 130331 193972 130332 194036
rect 130396 193972 130397 194036
rect 130331 193971 130397 193972
rect 128123 78436 128189 78437
rect 128123 78372 128124 78436
rect 128188 78372 128189 78436
rect 128123 78371 128189 78372
rect 126835 78300 126901 78301
rect 126835 78236 126836 78300
rect 126900 78236 126901 78300
rect 126835 78235 126901 78236
rect 126467 77620 126533 77621
rect 126467 77556 126468 77620
rect 126532 77556 126533 77620
rect 126467 77555 126533 77556
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 120579 31788 120645 31789
rect 120579 31724 120580 31788
rect 120644 31724 120645 31788
rect 120579 31723 120645 31724
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 130334 77485 130394 193971
rect 130518 81157 130578 197371
rect 130702 81293 130762 197507
rect 130699 81292 130765 81293
rect 130699 81228 130700 81292
rect 130764 81228 130765 81292
rect 130699 81227 130765 81228
rect 130515 81156 130581 81157
rect 130515 81092 130516 81156
rect 130580 81092 130581 81156
rect 130515 81091 130581 81092
rect 130886 78709 130946 198459
rect 133278 197709 133338 198690
rect 133459 198660 133525 198661
rect 133459 198596 133460 198660
rect 133524 198596 133525 198660
rect 133459 198595 133525 198596
rect 133275 197708 133341 197709
rect 133275 197644 133276 197708
rect 133340 197644 133341 197708
rect 133275 197643 133341 197644
rect 133091 196212 133157 196213
rect 133091 196148 133092 196212
rect 133156 196148 133157 196212
rect 133091 196147 133157 196148
rect 131619 196076 131685 196077
rect 131619 196012 131620 196076
rect 131684 196012 131685 196076
rect 131619 196011 131685 196012
rect 131622 79797 131682 196011
rect 131803 195940 131869 195941
rect 131803 195876 131804 195940
rect 131868 195876 131869 195940
rect 131803 195875 131869 195876
rect 131619 79796 131685 79797
rect 131619 79732 131620 79796
rect 131684 79732 131685 79796
rect 131619 79731 131685 79732
rect 130883 78708 130949 78709
rect 130883 78644 130884 78708
rect 130948 78644 130949 78708
rect 130883 78643 130949 78644
rect 131806 78029 131866 195875
rect 132171 195668 132237 195669
rect 132171 195604 132172 195668
rect 132236 195604 132237 195668
rect 132171 195603 132237 195604
rect 131987 139364 132053 139365
rect 131987 139300 131988 139364
rect 132052 139300 132053 139364
rect 131987 139299 132053 139300
rect 131990 79389 132050 139299
rect 132174 80613 132234 195603
rect 132171 80612 132237 80613
rect 132171 80548 132172 80612
rect 132236 80548 132237 80612
rect 132171 80547 132237 80548
rect 132907 79932 132973 79933
rect 132907 79868 132908 79932
rect 132972 79868 132973 79932
rect 132907 79867 132973 79868
rect 131987 79388 132053 79389
rect 131987 79324 131988 79388
rect 132052 79324 132053 79388
rect 131987 79323 132053 79324
rect 132910 78573 132970 79867
rect 133094 79797 133154 196147
rect 133275 196076 133341 196077
rect 133275 196012 133276 196076
rect 133340 196012 133341 196076
rect 133275 196011 133341 196012
rect 133091 79796 133157 79797
rect 133091 79732 133092 79796
rect 133156 79732 133157 79796
rect 133091 79731 133157 79732
rect 133278 79661 133338 196011
rect 133275 79660 133341 79661
rect 133275 79596 133276 79660
rect 133340 79596 133341 79660
rect 133275 79595 133341 79596
rect 133462 78573 133522 198595
rect 134379 197980 134445 197981
rect 134379 197916 134380 197980
rect 134444 197916 134445 197980
rect 134379 197915 134445 197916
rect 134563 197980 134629 197981
rect 134563 197916 134564 197980
rect 134628 197916 134629 197980
rect 134563 197915 134629 197916
rect 133643 197844 133709 197845
rect 133643 197780 133644 197844
rect 133708 197780 133709 197844
rect 133643 197779 133709 197780
rect 133646 79797 133706 197779
rect 134382 80069 134442 197915
rect 134566 81973 134626 197915
rect 134563 81972 134629 81973
rect 134563 81908 134564 81972
rect 134628 81908 134629 81972
rect 134563 81907 134629 81908
rect 134379 80068 134445 80069
rect 134379 80004 134380 80068
rect 134444 80004 134445 80068
rect 134379 80003 134445 80004
rect 133643 79796 133709 79797
rect 133643 79732 133644 79796
rect 133708 79732 133709 79796
rect 133643 79731 133709 79732
rect 132907 78572 132973 78573
rect 132907 78508 132908 78572
rect 132972 78508 132973 78572
rect 132907 78507 132973 78508
rect 133459 78572 133525 78573
rect 133459 78508 133460 78572
rect 133524 78508 133525 78572
rect 133459 78507 133525 78508
rect 131803 78028 131869 78029
rect 131803 77964 131804 78028
rect 131868 77964 131869 78028
rect 131803 77963 131869 77964
rect 130331 77484 130397 77485
rect 130331 77420 130332 77484
rect 130396 77420 130397 77484
rect 130331 77419 130397 77420
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 61954 132914 78000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 132294 25954 132914 61398
rect 133462 36549 133522 78507
rect 133646 66877 133706 79731
rect 134195 79660 134261 79661
rect 134195 79596 134196 79660
rect 134260 79596 134261 79660
rect 134195 79595 134261 79596
rect 134011 75988 134077 75989
rect 134011 75924 134012 75988
rect 134076 75924 134077 75988
rect 134011 75923 134077 75924
rect 133643 66876 133709 66877
rect 133643 66812 133644 66876
rect 133708 66812 133709 66876
rect 133643 66811 133709 66812
rect 134014 50965 134074 75923
rect 134198 52461 134258 79595
rect 134382 76669 134442 80003
rect 134563 79932 134629 79933
rect 134563 79868 134564 79932
rect 134628 79930 134629 79932
rect 134750 79930 134810 199819
rect 135851 199068 135917 199069
rect 135851 199004 135852 199068
rect 135916 199004 135917 199068
rect 135851 199003 135917 199004
rect 134931 197844 134997 197845
rect 134931 197780 134932 197844
rect 134996 197780 134997 197844
rect 134931 197779 134997 197780
rect 134628 79870 134810 79930
rect 134628 79868 134629 79870
rect 134563 79867 134629 79868
rect 134747 79796 134813 79797
rect 134747 79732 134748 79796
rect 134812 79732 134813 79796
rect 134747 79731 134813 79732
rect 134750 77349 134810 79731
rect 134934 79661 134994 197779
rect 135483 191044 135549 191045
rect 135483 190980 135484 191044
rect 135548 190980 135549 191044
rect 135483 190979 135549 190980
rect 135115 81972 135181 81973
rect 135115 81908 135116 81972
rect 135180 81908 135181 81972
rect 135115 81907 135181 81908
rect 135118 79797 135178 81907
rect 135115 79796 135181 79797
rect 135115 79732 135116 79796
rect 135180 79732 135181 79796
rect 135115 79731 135181 79732
rect 134931 79660 134997 79661
rect 134931 79596 134932 79660
rect 134996 79596 134997 79660
rect 134931 79595 134997 79596
rect 135486 78301 135546 190979
rect 135854 79933 135914 199003
rect 135851 79932 135917 79933
rect 135851 79868 135852 79932
rect 135916 79868 135917 79932
rect 135851 79867 135917 79868
rect 135854 78573 135914 79867
rect 135851 78572 135917 78573
rect 135851 78508 135852 78572
rect 135916 78508 135917 78572
rect 135851 78507 135917 78508
rect 135483 78300 135549 78301
rect 135483 78236 135484 78300
rect 135548 78236 135549 78300
rect 135483 78235 135549 78236
rect 136038 77893 136098 199819
rect 136403 199748 136469 199749
rect 136403 199684 136404 199748
rect 136468 199684 136469 199748
rect 136403 199683 136469 199684
rect 136406 199069 136466 199683
rect 136590 199613 136650 200499
rect 138059 200428 138125 200429
rect 138059 200364 138060 200428
rect 138124 200364 138125 200428
rect 138059 200363 138125 200364
rect 138062 200157 138122 200363
rect 138059 200156 138125 200157
rect 138059 200092 138060 200156
rect 138124 200092 138125 200156
rect 138059 200091 138125 200092
rect 138611 200020 138677 200021
rect 138611 199956 138612 200020
rect 138676 199956 138677 200020
rect 138611 199955 138677 199956
rect 137139 199748 137205 199749
rect 137139 199684 137140 199748
rect 137204 199684 137205 199748
rect 137139 199683 137205 199684
rect 137691 199748 137757 199749
rect 137691 199684 137692 199748
rect 137756 199684 137757 199748
rect 137691 199683 137757 199684
rect 136587 199612 136653 199613
rect 136587 199548 136588 199612
rect 136652 199548 136653 199612
rect 136587 199547 136653 199548
rect 136403 199068 136469 199069
rect 136403 199004 136404 199068
rect 136468 199004 136469 199068
rect 136403 199003 136469 199004
rect 136587 197844 136653 197845
rect 136587 197780 136588 197844
rect 136652 197780 136653 197844
rect 136587 197779 136653 197780
rect 136219 191180 136285 191181
rect 136219 191116 136220 191180
rect 136284 191116 136285 191180
rect 136219 191115 136285 191116
rect 136222 79661 136282 191115
rect 136590 79661 136650 197779
rect 137142 79933 137202 199683
rect 137507 197980 137573 197981
rect 137507 197916 137508 197980
rect 137572 197916 137573 197980
rect 137507 197915 137573 197916
rect 137323 81428 137389 81429
rect 137323 81364 137324 81428
rect 137388 81364 137389 81428
rect 137323 81363 137389 81364
rect 137139 79932 137205 79933
rect 137139 79868 137140 79932
rect 137204 79868 137205 79932
rect 137139 79867 137205 79868
rect 136955 79796 137021 79797
rect 136955 79732 136956 79796
rect 137020 79732 137021 79796
rect 136955 79731 137021 79732
rect 136219 79660 136285 79661
rect 136219 79596 136220 79660
rect 136284 79596 136285 79660
rect 136219 79595 136285 79596
rect 136587 79660 136653 79661
rect 136587 79596 136588 79660
rect 136652 79596 136653 79660
rect 136587 79595 136653 79596
rect 136958 78434 137018 79731
rect 137142 78573 137202 79867
rect 137326 79797 137386 81363
rect 137510 79933 137570 197915
rect 137694 79933 137754 199683
rect 138243 80340 138309 80341
rect 138243 80276 138244 80340
rect 138308 80276 138309 80340
rect 138243 80275 138309 80276
rect 137507 79932 137573 79933
rect 137507 79868 137508 79932
rect 137572 79868 137573 79932
rect 137507 79867 137573 79868
rect 137691 79932 137757 79933
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 137323 79796 137389 79797
rect 137323 79732 137324 79796
rect 137388 79732 137389 79796
rect 137323 79731 137389 79732
rect 138059 79116 138125 79117
rect 138059 79052 138060 79116
rect 138124 79114 138125 79116
rect 138246 79114 138306 80275
rect 138614 79661 138674 199955
rect 138795 199884 138861 199885
rect 138795 199820 138796 199884
rect 138860 199820 138861 199884
rect 138795 199819 138861 199820
rect 140635 199884 140701 199885
rect 140635 199820 140636 199884
rect 140700 199820 140701 199884
rect 140635 199819 140701 199820
rect 141003 199884 141069 199885
rect 141003 199820 141004 199884
rect 141068 199820 141069 199884
rect 141003 199819 141069 199820
rect 138798 79797 138858 199819
rect 140083 199748 140149 199749
rect 140083 199684 140084 199748
rect 140148 199684 140149 199748
rect 140083 199683 140149 199684
rect 139347 199612 139413 199613
rect 139347 199548 139348 199612
rect 139412 199548 139413 199612
rect 139347 199547 139413 199548
rect 139350 199069 139410 199547
rect 139347 199068 139413 199069
rect 139347 199004 139348 199068
rect 139412 199004 139413 199068
rect 139347 199003 139413 199004
rect 139163 198796 139229 198797
rect 139163 198732 139164 198796
rect 139228 198732 139229 198796
rect 139163 198731 139229 198732
rect 138979 183292 139045 183293
rect 138979 183228 138980 183292
rect 139044 183228 139045 183292
rect 138979 183227 139045 183228
rect 138982 79933 139042 183227
rect 138979 79932 139045 79933
rect 138979 79868 138980 79932
rect 139044 79868 139045 79932
rect 138979 79867 139045 79868
rect 138795 79796 138861 79797
rect 138795 79732 138796 79796
rect 138860 79732 138861 79796
rect 138795 79731 138861 79732
rect 139166 79661 139226 198731
rect 140086 198117 140146 199683
rect 140267 199068 140333 199069
rect 140267 199004 140268 199068
rect 140332 199004 140333 199068
rect 140267 199003 140333 199004
rect 139347 198116 139413 198117
rect 139347 198052 139348 198116
rect 139412 198052 139413 198116
rect 139347 198051 139413 198052
rect 140083 198116 140149 198117
rect 140083 198052 140084 198116
rect 140148 198052 140149 198116
rect 140083 198051 140149 198052
rect 139350 81565 139410 198051
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 139347 81564 139413 81565
rect 139347 81500 139348 81564
rect 139412 81500 139413 81564
rect 139347 81499 139413 81500
rect 139350 79797 139410 81499
rect 139531 79932 139597 79933
rect 139531 79868 139532 79932
rect 139596 79868 139597 79932
rect 139531 79867 139597 79868
rect 139347 79796 139413 79797
rect 139347 79732 139348 79796
rect 139412 79732 139413 79796
rect 139347 79731 139413 79732
rect 138427 79660 138493 79661
rect 138427 79596 138428 79660
rect 138492 79596 138493 79660
rect 138427 79595 138493 79596
rect 138611 79660 138677 79661
rect 138611 79596 138612 79660
rect 138676 79596 138677 79660
rect 138611 79595 138677 79596
rect 139163 79660 139229 79661
rect 139163 79596 139164 79660
rect 139228 79596 139229 79660
rect 139163 79595 139229 79596
rect 138124 79054 138306 79114
rect 138124 79052 138125 79054
rect 138059 79051 138125 79052
rect 137139 78572 137205 78573
rect 137139 78508 137140 78572
rect 137204 78508 137205 78572
rect 137139 78507 137205 78508
rect 138059 78572 138125 78573
rect 138059 78508 138060 78572
rect 138124 78508 138125 78572
rect 138059 78507 138125 78508
rect 136958 78374 137754 78434
rect 136035 77892 136101 77893
rect 136035 77828 136036 77892
rect 136100 77828 136101 77892
rect 136035 77827 136101 77828
rect 134747 77348 134813 77349
rect 134747 77284 134748 77348
rect 134812 77284 134813 77348
rect 134747 77283 134813 77284
rect 134931 77212 134997 77213
rect 134931 77148 134932 77212
rect 134996 77148 134997 77212
rect 134931 77147 134997 77148
rect 134379 76668 134445 76669
rect 134379 76604 134380 76668
rect 134444 76604 134445 76668
rect 134379 76603 134445 76604
rect 134379 74220 134445 74221
rect 134379 74156 134380 74220
rect 134444 74156 134445 74220
rect 134379 74155 134445 74156
rect 134382 57901 134442 74155
rect 134379 57900 134445 57901
rect 134379 57836 134380 57900
rect 134444 57836 134445 57900
rect 134379 57835 134445 57836
rect 134195 52460 134261 52461
rect 134195 52396 134196 52460
rect 134260 52396 134261 52460
rect 134195 52395 134261 52396
rect 134011 50964 134077 50965
rect 134011 50900 134012 50964
rect 134076 50900 134077 50964
rect 134011 50899 134077 50900
rect 133459 36548 133525 36549
rect 133459 36484 133460 36548
rect 133524 36484 133525 36548
rect 133459 36483 133525 36484
rect 134934 33829 134994 77147
rect 135667 75988 135733 75989
rect 135667 75924 135668 75988
rect 135732 75924 135733 75988
rect 135667 75923 135733 75924
rect 135851 75988 135917 75989
rect 135851 75924 135852 75988
rect 135916 75924 135917 75988
rect 135851 75923 135917 75924
rect 135483 75852 135549 75853
rect 135483 75788 135484 75852
rect 135548 75788 135549 75852
rect 135483 75787 135549 75788
rect 135486 49605 135546 75787
rect 135670 67557 135730 75923
rect 135667 67556 135733 67557
rect 135667 67492 135668 67556
rect 135732 67492 135733 67556
rect 135667 67491 135733 67492
rect 135483 49604 135549 49605
rect 135483 49540 135484 49604
rect 135548 49540 135549 49604
rect 135483 49539 135549 49540
rect 135854 48245 135914 75923
rect 136794 66454 137414 78000
rect 137507 74900 137573 74901
rect 137507 74836 137508 74900
rect 137572 74836 137573 74900
rect 137507 74835 137573 74836
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 137510 66197 137570 74835
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 137507 66196 137573 66197
rect 137507 66132 137508 66196
rect 137572 66132 137573 66196
rect 137507 66131 137573 66132
rect 135851 48244 135917 48245
rect 135851 48180 135852 48244
rect 135916 48180 135917 48244
rect 135851 48179 135917 48180
rect 134931 33828 134997 33829
rect 134931 33764 134932 33828
rect 134996 33764 134997 33828
rect 134931 33763 134997 33764
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 65898
rect 137694 46885 137754 78374
rect 137691 46884 137757 46885
rect 137691 46820 137692 46884
rect 137756 46820 137757 46884
rect 137691 46819 137757 46820
rect 138062 44165 138122 78507
rect 138243 77620 138309 77621
rect 138243 77556 138244 77620
rect 138308 77556 138309 77620
rect 138243 77555 138309 77556
rect 138246 55181 138306 77555
rect 138430 57765 138490 79595
rect 138611 77756 138677 77757
rect 138611 77692 138612 77756
rect 138676 77692 138677 77756
rect 138611 77691 138677 77692
rect 138614 63477 138674 77691
rect 139166 77485 139226 79595
rect 139347 78708 139413 78709
rect 139347 78644 139348 78708
rect 139412 78644 139413 78708
rect 139347 78643 139413 78644
rect 139163 77484 139229 77485
rect 139163 77420 139164 77484
rect 139228 77420 139229 77484
rect 139163 77419 139229 77420
rect 139350 75717 139410 78643
rect 139347 75716 139413 75717
rect 139347 75652 139348 75716
rect 139412 75652 139413 75716
rect 139347 75651 139413 75652
rect 139534 72997 139594 79867
rect 140270 79797 140330 199003
rect 140451 198116 140517 198117
rect 140451 198052 140452 198116
rect 140516 198052 140517 198116
rect 140451 198051 140517 198052
rect 140267 79796 140333 79797
rect 140267 79732 140268 79796
rect 140332 79732 140333 79796
rect 140267 79731 140333 79732
rect 139715 79660 139781 79661
rect 139715 79596 139716 79660
rect 139780 79596 139781 79660
rect 139715 79595 139781 79596
rect 139718 74085 139778 79595
rect 140270 77349 140330 79731
rect 140454 78981 140514 198051
rect 140638 79661 140698 199819
rect 140819 199748 140885 199749
rect 140819 199684 140820 199748
rect 140884 199684 140885 199748
rect 140819 199683 140885 199684
rect 140822 197029 140882 199683
rect 141006 197981 141066 199819
rect 141558 199613 141618 200635
rect 150203 200292 150269 200293
rect 150203 200228 150204 200292
rect 150268 200228 150269 200292
rect 150203 200227 150269 200228
rect 170259 200292 170325 200293
rect 170259 200228 170260 200292
rect 170324 200228 170325 200292
rect 170259 200227 170325 200228
rect 150019 200156 150085 200157
rect 150019 200092 150020 200156
rect 150084 200092 150085 200156
rect 150019 200091 150085 200092
rect 142475 199884 142541 199885
rect 142475 199820 142476 199884
rect 142540 199820 142541 199884
rect 142475 199819 142541 199820
rect 144499 199884 144565 199885
rect 144499 199820 144500 199884
rect 144564 199820 144565 199884
rect 144499 199819 144565 199820
rect 145419 199884 145485 199885
rect 145419 199820 145420 199884
rect 145484 199820 145485 199884
rect 145419 199819 145485 199820
rect 147075 199884 147141 199885
rect 147075 199820 147076 199884
rect 147140 199820 147141 199884
rect 147075 199819 147141 199820
rect 147811 199884 147877 199885
rect 147811 199820 147812 199884
rect 147876 199820 147877 199884
rect 147811 199819 147877 199820
rect 147995 199884 148061 199885
rect 147995 199820 147996 199884
rect 148060 199820 148061 199884
rect 147995 199819 148061 199820
rect 148547 199884 148613 199885
rect 148547 199820 148548 199884
rect 148612 199820 148613 199884
rect 148547 199819 148613 199820
rect 149651 199884 149717 199885
rect 149651 199820 149652 199884
rect 149716 199820 149717 199884
rect 149651 199819 149717 199820
rect 141555 199612 141621 199613
rect 141555 199548 141556 199612
rect 141620 199548 141621 199612
rect 141555 199547 141621 199548
rect 141003 197980 141069 197981
rect 141003 197916 141004 197980
rect 141068 197916 141069 197980
rect 141003 197915 141069 197916
rect 140819 197028 140885 197029
rect 140819 196964 140820 197028
rect 140884 196964 140885 197028
rect 140819 196963 140885 196964
rect 140819 196076 140885 196077
rect 140819 196012 140820 196076
rect 140884 196012 140885 196076
rect 140819 196011 140885 196012
rect 140635 79660 140701 79661
rect 140635 79596 140636 79660
rect 140700 79596 140701 79660
rect 140635 79595 140701 79596
rect 140451 78980 140517 78981
rect 140451 78916 140452 78980
rect 140516 78916 140517 78980
rect 140451 78915 140517 78916
rect 140638 77757 140698 79595
rect 140635 77756 140701 77757
rect 140635 77692 140636 77756
rect 140700 77692 140701 77756
rect 140635 77691 140701 77692
rect 140822 77485 140882 196011
rect 141003 188868 141069 188869
rect 141003 188804 141004 188868
rect 141068 188804 141069 188868
rect 141003 188803 141069 188804
rect 141006 79933 141066 188803
rect 141294 178954 141914 198000
rect 142478 196485 142538 199819
rect 144131 198116 144197 198117
rect 144131 198052 144132 198116
rect 144196 198052 144197 198116
rect 144131 198051 144197 198052
rect 142659 197980 142725 197981
rect 142659 197916 142660 197980
rect 142724 197916 142725 197980
rect 142659 197915 142725 197916
rect 142475 196484 142541 196485
rect 142475 196420 142476 196484
rect 142540 196420 142541 196484
rect 142475 196419 142541 196420
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 142475 149700 142541 149701
rect 142475 149636 142476 149700
rect 142540 149636 142541 149700
rect 142475 149635 142541 149636
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 141371 141268 141437 141269
rect 141371 141204 141372 141268
rect 141436 141204 141437 141268
rect 141371 141203 141437 141204
rect 141003 79932 141069 79933
rect 141003 79868 141004 79932
rect 141068 79868 141069 79932
rect 141003 79867 141069 79868
rect 141003 79796 141069 79797
rect 141003 79732 141004 79796
rect 141068 79732 141069 79796
rect 141003 79731 141069 79732
rect 140819 77484 140885 77485
rect 140819 77420 140820 77484
rect 140884 77420 140885 77484
rect 140819 77419 140885 77420
rect 140267 77348 140333 77349
rect 140267 77284 140268 77348
rect 140332 77284 140333 77348
rect 140267 77283 140333 77284
rect 140819 77348 140885 77349
rect 140819 77284 140820 77348
rect 140884 77284 140885 77348
rect 140819 77283 140885 77284
rect 139715 74084 139781 74085
rect 139715 74020 139716 74084
rect 139780 74020 139781 74084
rect 139715 74019 139781 74020
rect 140822 73949 140882 77283
rect 141006 75581 141066 79731
rect 141374 79661 141434 141203
rect 141555 141132 141621 141133
rect 141555 141068 141556 141132
rect 141620 141068 141621 141132
rect 141555 141067 141621 141068
rect 141558 79797 141618 141067
rect 141555 79796 141621 79797
rect 141555 79732 141556 79796
rect 141620 79732 141621 79796
rect 141555 79731 141621 79732
rect 141371 79660 141437 79661
rect 141371 79596 141372 79660
rect 141436 79596 141437 79660
rect 141371 79595 141437 79596
rect 142107 78980 142173 78981
rect 142107 78916 142108 78980
rect 142172 78916 142173 78980
rect 142107 78915 142173 78916
rect 141003 75580 141069 75581
rect 141003 75516 141004 75580
rect 141068 75516 141069 75580
rect 141003 75515 141069 75516
rect 140819 73948 140885 73949
rect 140819 73884 140820 73948
rect 140884 73884 140885 73948
rect 140819 73883 140885 73884
rect 139531 72996 139597 72997
rect 139531 72932 139532 72996
rect 139596 72932 139597 72996
rect 139531 72931 139597 72932
rect 141294 70954 141914 78000
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 142110 70413 142170 78915
rect 142478 78437 142538 149635
rect 142662 78981 142722 197915
rect 143579 197028 143645 197029
rect 143579 196964 143580 197028
rect 143644 196964 143645 197028
rect 143579 196963 143645 196964
rect 142843 195396 142909 195397
rect 142843 195332 142844 195396
rect 142908 195332 142909 195396
rect 142843 195331 142909 195332
rect 142846 81429 142906 195331
rect 143582 189685 143642 196963
rect 143579 189684 143645 189685
rect 143579 189620 143580 189684
rect 143644 189620 143645 189684
rect 143579 189619 143645 189620
rect 144134 144669 144194 198051
rect 144502 193221 144562 199819
rect 145422 199069 145482 199819
rect 145603 199748 145669 199749
rect 145603 199684 145604 199748
rect 145668 199684 145669 199748
rect 145603 199683 145669 199684
rect 145419 199068 145485 199069
rect 145419 199004 145420 199068
rect 145484 199004 145485 199068
rect 145419 199003 145485 199004
rect 145606 198522 145666 199683
rect 146891 198932 146957 198933
rect 146891 198868 146892 198932
rect 146956 198868 146957 198932
rect 146891 198867 146957 198868
rect 145422 198462 145666 198522
rect 144683 197980 144749 197981
rect 144683 197916 144684 197980
rect 144748 197916 144749 197980
rect 144683 197915 144749 197916
rect 144686 195397 144746 197915
rect 145235 196076 145301 196077
rect 145235 196012 145236 196076
rect 145300 196012 145301 196076
rect 145235 196011 145301 196012
rect 144683 195396 144749 195397
rect 144683 195332 144684 195396
rect 144748 195332 144749 195396
rect 144683 195331 144749 195332
rect 144499 193220 144565 193221
rect 144499 193156 144500 193220
rect 144564 193156 144565 193220
rect 144499 193155 144565 193156
rect 144131 144668 144197 144669
rect 144131 144604 144132 144668
rect 144196 144604 144197 144668
rect 144131 144603 144197 144604
rect 142843 81428 142909 81429
rect 142843 81364 142844 81428
rect 142908 81364 142909 81428
rect 142843 81363 142909 81364
rect 143211 81292 143277 81293
rect 143211 81228 143212 81292
rect 143276 81228 143277 81292
rect 143211 81227 143277 81228
rect 143027 79932 143093 79933
rect 143027 79868 143028 79932
rect 143092 79868 143093 79932
rect 143027 79867 143093 79868
rect 142659 78980 142725 78981
rect 142659 78916 142660 78980
rect 142724 78916 142725 78980
rect 142659 78915 142725 78916
rect 142475 78436 142541 78437
rect 142475 78372 142476 78436
rect 142540 78372 142541 78436
rect 142475 78371 142541 78372
rect 143030 77213 143090 79867
rect 143214 78981 143274 81227
rect 143395 81156 143461 81157
rect 143395 81092 143396 81156
rect 143460 81092 143461 81156
rect 143395 81091 143461 81092
rect 143211 78980 143277 78981
rect 143211 78916 143212 78980
rect 143276 78916 143277 78980
rect 143211 78915 143277 78916
rect 143398 78709 143458 81091
rect 144867 80884 144933 80885
rect 144867 80820 144868 80884
rect 144932 80820 144933 80884
rect 144867 80819 144933 80820
rect 144315 79932 144381 79933
rect 144315 79868 144316 79932
rect 144380 79868 144381 79932
rect 144315 79867 144381 79868
rect 143395 78708 143461 78709
rect 143395 78644 143396 78708
rect 143460 78644 143461 78708
rect 143395 78643 143461 78644
rect 143027 77212 143093 77213
rect 143027 77148 143028 77212
rect 143092 77148 143093 77212
rect 143027 77147 143093 77148
rect 144131 71092 144197 71093
rect 144131 71028 144132 71092
rect 144196 71028 144197 71092
rect 144131 71027 144197 71028
rect 138611 63476 138677 63477
rect 138611 63412 138612 63476
rect 138676 63412 138677 63476
rect 138611 63411 138677 63412
rect 138427 57764 138493 57765
rect 138427 57700 138428 57764
rect 138492 57700 138493 57764
rect 138427 57699 138493 57700
rect 138243 55180 138309 55181
rect 138243 55116 138244 55180
rect 138308 55116 138309 55180
rect 138243 55115 138309 55116
rect 138059 44164 138125 44165
rect 138059 44100 138060 44164
rect 138124 44100 138125 44164
rect 138059 44099 138125 44100
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 70398
rect 142107 70412 142173 70413
rect 142107 70348 142108 70412
rect 142172 70348 142173 70412
rect 142107 70347 142173 70348
rect 142107 64972 142173 64973
rect 142107 64908 142108 64972
rect 142172 64908 142173 64972
rect 142107 64907 142173 64908
rect 142110 64701 142170 64907
rect 142107 64700 142173 64701
rect 142107 64636 142108 64700
rect 142172 64636 142173 64700
rect 142107 64635 142173 64636
rect 142107 55316 142173 55317
rect 142107 55252 142108 55316
rect 142172 55252 142173 55316
rect 142107 55251 142173 55252
rect 142110 55045 142170 55251
rect 142107 55044 142173 55045
rect 142107 54980 142108 55044
rect 142172 54980 142173 55044
rect 142107 54979 142173 54980
rect 142107 45660 142173 45661
rect 142107 45596 142108 45660
rect 142172 45596 142173 45660
rect 142107 45595 142173 45596
rect 142110 45525 142170 45595
rect 142107 45524 142173 45525
rect 142107 45460 142108 45524
rect 142172 45460 142173 45524
rect 142107 45459 142173 45460
rect 142107 36140 142173 36141
rect 142107 36076 142108 36140
rect 142172 36076 142173 36140
rect 142107 36075 142173 36076
rect 142110 35910 142170 36075
rect 142110 35869 142354 35910
rect 142110 35868 142357 35869
rect 142110 35850 142292 35868
rect 142291 35804 142292 35850
rect 142356 35804 142357 35868
rect 142291 35803 142357 35804
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 142107 26348 142173 26349
rect 142107 26284 142108 26348
rect 142172 26284 142173 26348
rect 142107 26283 142173 26284
rect 142110 26213 142170 26283
rect 142107 26212 142173 26213
rect 142107 26148 142108 26212
rect 142172 26148 142173 26212
rect 142107 26147 142173 26148
rect 142291 16692 142357 16693
rect 142291 16690 142292 16692
rect 142110 16630 142292 16690
rect 142110 16421 142170 16630
rect 142291 16628 142292 16630
rect 142356 16628 142357 16692
rect 142291 16627 142357 16628
rect 142107 16420 142173 16421
rect 142107 16356 142108 16420
rect 142172 16356 142173 16420
rect 142107 16355 142173 16356
rect 142107 7036 142173 7037
rect 142107 6972 142108 7036
rect 142172 6972 142173 7036
rect 142107 6971 142173 6972
rect 142110 6901 142170 6971
rect 142107 6900 142173 6901
rect 142107 6836 142108 6900
rect 142172 6836 142173 6900
rect 142107 6835 142173 6836
rect 144134 4861 144194 71027
rect 144318 68645 144378 79867
rect 144870 79797 144930 80819
rect 145051 80476 145117 80477
rect 145051 80412 145052 80476
rect 145116 80412 145117 80476
rect 145051 80411 145117 80412
rect 145054 79933 145114 80411
rect 145051 79932 145117 79933
rect 145051 79868 145052 79932
rect 145116 79868 145117 79932
rect 145051 79867 145117 79868
rect 144499 79796 144565 79797
rect 144499 79732 144500 79796
rect 144564 79732 144565 79796
rect 144499 79731 144565 79732
rect 144867 79796 144933 79797
rect 144867 79732 144868 79796
rect 144932 79732 144933 79796
rect 144867 79731 144933 79732
rect 144502 70005 144562 79731
rect 145238 79253 145298 196011
rect 145422 80069 145482 198462
rect 145603 198252 145669 198253
rect 145603 198188 145604 198252
rect 145668 198188 145669 198252
rect 145603 198187 145669 198188
rect 145419 80068 145485 80069
rect 145419 80004 145420 80068
rect 145484 80004 145485 80068
rect 145419 80003 145485 80004
rect 145419 79932 145485 79933
rect 145419 79868 145420 79932
rect 145484 79868 145485 79932
rect 145419 79867 145485 79868
rect 145235 79252 145301 79253
rect 145235 79188 145236 79252
rect 145300 79188 145301 79252
rect 145235 79187 145301 79188
rect 145422 79117 145482 79867
rect 145419 79116 145485 79117
rect 145419 79052 145420 79116
rect 145484 79052 145485 79116
rect 145419 79051 145485 79052
rect 144683 74764 144749 74765
rect 144683 74700 144684 74764
rect 144748 74700 144749 74764
rect 144683 74699 144749 74700
rect 144499 70004 144565 70005
rect 144499 69940 144500 70004
rect 144564 69940 144565 70004
rect 144499 69939 144565 69940
rect 144315 68644 144381 68645
rect 144315 68580 144316 68644
rect 144380 68580 144381 68644
rect 144315 68579 144381 68580
rect 144318 15877 144378 68579
rect 144502 21317 144562 69939
rect 144686 68917 144746 74699
rect 145051 73948 145117 73949
rect 145051 73884 145052 73948
rect 145116 73884 145117 73948
rect 145051 73883 145117 73884
rect 145054 71365 145114 73883
rect 145422 72317 145482 79051
rect 145606 78981 145666 198187
rect 145794 183454 146414 198000
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 146894 79661 146954 198867
rect 146891 79660 146957 79661
rect 146891 79596 146892 79660
rect 146956 79596 146957 79660
rect 146891 79595 146957 79596
rect 147078 79117 147138 199819
rect 147814 196077 147874 199819
rect 147998 198933 148058 199819
rect 147995 198932 148061 198933
rect 147995 198868 147996 198932
rect 148060 198868 148061 198932
rect 147995 198867 148061 198868
rect 147811 196076 147877 196077
rect 147811 196012 147812 196076
rect 147876 196012 147877 196076
rect 147811 196011 147877 196012
rect 148550 195941 148610 199819
rect 148731 199748 148797 199749
rect 148731 199684 148732 199748
rect 148796 199684 148797 199748
rect 148731 199683 148797 199684
rect 148734 198933 148794 199683
rect 149654 199477 149714 199819
rect 149651 199476 149717 199477
rect 149651 199412 149652 199476
rect 149716 199412 149717 199476
rect 149651 199411 149717 199412
rect 148731 198932 148797 198933
rect 148731 198868 148732 198932
rect 148796 198868 148797 198932
rect 148731 198867 148797 198868
rect 148915 198660 148981 198661
rect 148915 198596 148916 198660
rect 148980 198596 148981 198660
rect 148915 198595 148981 198596
rect 148731 197572 148797 197573
rect 148731 197508 148732 197572
rect 148796 197508 148797 197572
rect 148731 197507 148797 197508
rect 148547 195940 148613 195941
rect 148547 195876 148548 195940
rect 148612 195876 148613 195940
rect 148547 195875 148613 195876
rect 147259 195532 147325 195533
rect 147259 195468 147260 195532
rect 147324 195468 147325 195532
rect 147259 195467 147325 195468
rect 147262 93870 147322 195467
rect 148179 191180 148245 191181
rect 148179 191116 148180 191180
rect 148244 191116 148245 191180
rect 148179 191115 148245 191116
rect 147262 93810 147506 93870
rect 146707 79116 146773 79117
rect 146707 79052 146708 79116
rect 146772 79052 146773 79116
rect 146707 79051 146773 79052
rect 147075 79116 147141 79117
rect 147075 79052 147076 79116
rect 147140 79052 147141 79116
rect 147075 79051 147141 79052
rect 145603 78980 145669 78981
rect 145603 78916 145604 78980
rect 145668 78916 145669 78980
rect 145603 78915 145669 78916
rect 145794 75454 146414 78000
rect 145603 75444 145669 75445
rect 145603 75380 145604 75444
rect 145668 75380 145669 75444
rect 145603 75379 145669 75380
rect 145419 72316 145485 72317
rect 145419 72252 145420 72316
rect 145484 72252 145485 72316
rect 145419 72251 145485 72252
rect 145051 71364 145117 71365
rect 145051 71300 145052 71364
rect 145116 71300 145117 71364
rect 145051 71299 145117 71300
rect 144683 68916 144749 68917
rect 144683 68852 144684 68916
rect 144748 68852 144749 68916
rect 144683 68851 144749 68852
rect 144686 50693 144746 68851
rect 145054 64890 145114 71299
rect 145606 68917 145666 75379
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145603 68916 145669 68917
rect 145603 68852 145604 68916
rect 145668 68852 145669 68916
rect 145603 68851 145669 68852
rect 145054 64830 145482 64890
rect 144683 50692 144749 50693
rect 144683 50628 144684 50692
rect 144748 50628 144749 50692
rect 144683 50627 144749 50628
rect 145422 27029 145482 64830
rect 145794 39454 146414 74898
rect 146710 44981 146770 79051
rect 147446 78029 147506 93810
rect 147995 81020 148061 81021
rect 147995 80956 147996 81020
rect 148060 80956 148061 81020
rect 147995 80955 148061 80956
rect 147998 79797 148058 80955
rect 147995 79796 148061 79797
rect 147995 79732 147996 79796
rect 148060 79732 148061 79796
rect 147995 79731 148061 79732
rect 148182 79658 148242 191115
rect 148363 191044 148429 191045
rect 148363 190980 148364 191044
rect 148428 190980 148429 191044
rect 148363 190979 148429 190980
rect 148366 79797 148426 190979
rect 148593 79932 148659 79933
rect 148593 79930 148594 79932
rect 148550 79868 148594 79930
rect 148658 79868 148659 79932
rect 148550 79867 148659 79868
rect 148363 79796 148429 79797
rect 148363 79732 148364 79796
rect 148428 79732 148429 79796
rect 148363 79731 148429 79732
rect 148550 79658 148610 79867
rect 148182 79598 148610 79658
rect 148179 79116 148245 79117
rect 148179 79052 148180 79116
rect 148244 79052 148245 79116
rect 148179 79051 148245 79052
rect 147443 78028 147509 78029
rect 147443 77964 147444 78028
rect 147508 77964 147509 78028
rect 147443 77963 147509 77964
rect 146891 77076 146957 77077
rect 146891 77012 146892 77076
rect 146956 77012 146957 77076
rect 146891 77011 146957 77012
rect 146894 66877 146954 77011
rect 148182 76805 148242 79051
rect 148363 78300 148429 78301
rect 148363 78236 148364 78300
rect 148428 78236 148429 78300
rect 148363 78235 148429 78236
rect 148179 76804 148245 76805
rect 148179 76740 148180 76804
rect 148244 76740 148245 76804
rect 148179 76739 148245 76740
rect 148182 67149 148242 76739
rect 148366 75037 148426 78235
rect 148550 77757 148610 79598
rect 148734 79253 148794 197507
rect 148731 79252 148797 79253
rect 148731 79188 148732 79252
rect 148796 79188 148797 79252
rect 148731 79187 148797 79188
rect 148918 78845 148978 198595
rect 149835 197028 149901 197029
rect 149835 196964 149836 197028
rect 149900 196964 149901 197028
rect 149835 196963 149901 196964
rect 149467 196892 149533 196893
rect 149467 196828 149468 196892
rect 149532 196828 149533 196892
rect 149467 196827 149533 196828
rect 149099 79796 149165 79797
rect 149099 79732 149100 79796
rect 149164 79732 149165 79796
rect 149099 79731 149165 79732
rect 148915 78844 148981 78845
rect 148915 78780 148916 78844
rect 148980 78780 148981 78844
rect 148915 78779 148981 78780
rect 149102 78706 149162 79731
rect 148918 78646 149162 78706
rect 148547 77756 148613 77757
rect 148547 77692 148548 77756
rect 148612 77692 148613 77756
rect 148547 77691 148613 77692
rect 148731 75988 148797 75989
rect 148731 75924 148732 75988
rect 148796 75924 148797 75988
rect 148731 75923 148797 75924
rect 148363 75036 148429 75037
rect 148363 74972 148364 75036
rect 148428 74972 148429 75036
rect 148363 74971 148429 74972
rect 148366 70410 148426 74971
rect 148366 70350 148610 70410
rect 148550 68373 148610 70350
rect 148734 70141 148794 75923
rect 148731 70140 148797 70141
rect 148731 70076 148732 70140
rect 148796 70076 148797 70140
rect 148731 70075 148797 70076
rect 148547 68372 148613 68373
rect 148547 68308 148548 68372
rect 148612 68308 148613 68372
rect 148547 68307 148613 68308
rect 148179 67148 148245 67149
rect 148179 67084 148180 67148
rect 148244 67084 148245 67148
rect 148179 67083 148245 67084
rect 146891 66876 146957 66877
rect 146891 66812 146892 66876
rect 146956 66812 146957 66876
rect 146891 66811 146957 66812
rect 146707 44980 146773 44981
rect 146707 44916 146708 44980
rect 146772 44916 146773 44980
rect 146707 44915 146773 44916
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145419 27028 145485 27029
rect 145419 26964 145420 27028
rect 145484 26964 145485 27028
rect 145419 26963 145485 26964
rect 144499 21316 144565 21317
rect 144499 21252 144500 21316
rect 144564 21252 144565 21316
rect 144499 21251 144565 21252
rect 144315 15876 144381 15877
rect 144315 15812 144316 15876
rect 144380 15812 144381 15876
rect 144315 15811 144381 15812
rect 144131 4860 144197 4861
rect 144131 4796 144132 4860
rect 144196 4796 144197 4860
rect 144131 4795 144197 4796
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3454 146414 38898
rect 148918 32469 148978 78646
rect 149099 78300 149165 78301
rect 149099 78236 149100 78300
rect 149164 78236 149165 78300
rect 149099 78235 149165 78236
rect 149102 72725 149162 78235
rect 149470 77757 149530 196827
rect 149651 196484 149717 196485
rect 149651 196420 149652 196484
rect 149716 196420 149717 196484
rect 149651 196419 149717 196420
rect 149654 79797 149714 196419
rect 149651 79796 149717 79797
rect 149651 79732 149652 79796
rect 149716 79732 149717 79796
rect 149651 79731 149717 79732
rect 149467 77756 149533 77757
rect 149467 77692 149468 77756
rect 149532 77692 149533 77756
rect 149467 77691 149533 77692
rect 149654 75930 149714 79731
rect 149838 79661 149898 196963
rect 149835 79660 149901 79661
rect 149835 79596 149836 79660
rect 149900 79596 149901 79660
rect 149835 79595 149901 79596
rect 149838 79117 149898 79595
rect 150022 79117 150082 200091
rect 150206 199477 150266 200227
rect 151307 200020 151373 200021
rect 151307 199956 151308 200020
rect 151372 199956 151373 200020
rect 151307 199955 151373 199956
rect 151491 200020 151557 200021
rect 151491 199956 151492 200020
rect 151556 199956 151557 200020
rect 151491 199955 151557 199956
rect 153515 200020 153581 200021
rect 153515 199956 153516 200020
rect 153580 199956 153581 200020
rect 153515 199955 153581 199956
rect 165291 200020 165357 200021
rect 165291 199956 165292 200020
rect 165356 199956 165357 200020
rect 165291 199955 165357 199956
rect 168787 200020 168853 200021
rect 168787 199956 168788 200020
rect 168852 199956 168853 200020
rect 168787 199955 168853 199956
rect 150387 199884 150453 199885
rect 150387 199820 150388 199884
rect 150452 199820 150453 199884
rect 150387 199819 150453 199820
rect 150755 199884 150821 199885
rect 150755 199820 150756 199884
rect 150820 199820 150821 199884
rect 150755 199819 150821 199820
rect 150203 199476 150269 199477
rect 150203 199412 150204 199476
rect 150268 199412 150269 199476
rect 150203 199411 150269 199412
rect 150390 198525 150450 199819
rect 150758 198797 150818 199819
rect 150755 198796 150821 198797
rect 150755 198732 150756 198796
rect 150820 198732 150821 198796
rect 150755 198731 150821 198732
rect 150387 198524 150453 198525
rect 150387 198460 150388 198524
rect 150452 198460 150453 198524
rect 150387 198459 150453 198460
rect 150294 187954 150914 198000
rect 151310 197029 151370 199955
rect 151307 197028 151373 197029
rect 151307 196964 151308 197028
rect 151372 196964 151373 197028
rect 151307 196963 151373 196964
rect 151494 196210 151554 199955
rect 152043 199884 152109 199885
rect 152043 199820 152044 199884
rect 152108 199820 152109 199884
rect 152043 199819 152109 199820
rect 152227 199884 152293 199885
rect 152227 199820 152228 199884
rect 152292 199820 152293 199884
rect 152779 199884 152845 199885
rect 152779 199882 152780 199884
rect 152227 199819 152293 199820
rect 152598 199822 152780 199882
rect 152046 199477 152106 199819
rect 151675 199476 151741 199477
rect 151675 199412 151676 199476
rect 151740 199412 151741 199476
rect 151675 199411 151741 199412
rect 152043 199476 152109 199477
rect 152043 199412 152044 199476
rect 152108 199412 152109 199476
rect 152043 199411 152109 199412
rect 151678 196757 151738 199411
rect 151675 196756 151741 196757
rect 151675 196692 151676 196756
rect 151740 196692 151741 196756
rect 151675 196691 151741 196692
rect 151310 196150 151554 196210
rect 151123 195668 151189 195669
rect 151123 195604 151124 195668
rect 151188 195604 151189 195668
rect 151123 195603 151189 195604
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 142000 150914 151398
rect 150755 139364 150821 139365
rect 150755 139300 150756 139364
rect 150820 139300 150821 139364
rect 150755 139299 150821 139300
rect 150758 80205 150818 139299
rect 151126 85590 151186 195603
rect 150942 85530 151186 85590
rect 150755 80204 150821 80205
rect 150755 80140 150756 80204
rect 150820 80140 150821 80204
rect 150755 80139 150821 80140
rect 150203 79932 150269 79933
rect 150203 79868 150204 79932
rect 150268 79868 150269 79932
rect 150203 79867 150269 79868
rect 150387 79932 150453 79933
rect 150387 79868 150388 79932
rect 150452 79868 150453 79932
rect 150387 79867 150453 79868
rect 149835 79116 149901 79117
rect 149835 79052 149836 79116
rect 149900 79052 149901 79116
rect 149835 79051 149901 79052
rect 150019 79116 150085 79117
rect 150019 79052 150020 79116
rect 150084 79052 150085 79116
rect 150019 79051 150085 79052
rect 150206 78434 150266 79867
rect 149286 75870 149714 75930
rect 149838 78374 150266 78434
rect 149099 72724 149165 72725
rect 149099 72660 149100 72724
rect 149164 72660 149165 72724
rect 149099 72659 149165 72660
rect 149286 42125 149346 75870
rect 149838 73810 149898 78374
rect 150390 78162 150450 79867
rect 150758 78437 150818 80139
rect 150942 79933 151002 85530
rect 150939 79932 151005 79933
rect 150939 79868 150940 79932
rect 151004 79868 151005 79932
rect 150939 79867 151005 79868
rect 151310 79661 151370 196150
rect 151491 196076 151557 196077
rect 151491 196012 151492 196076
rect 151556 196012 151557 196076
rect 151491 196011 151557 196012
rect 151494 79933 151554 196011
rect 152230 79933 152290 199819
rect 152411 183564 152477 183565
rect 152411 183500 152412 183564
rect 152476 183500 152477 183564
rect 152411 183499 152477 183500
rect 151491 79932 151557 79933
rect 151491 79868 151492 79932
rect 151556 79868 151557 79932
rect 151491 79867 151557 79868
rect 152227 79932 152293 79933
rect 152227 79868 152228 79932
rect 152292 79868 152293 79932
rect 152227 79867 152293 79868
rect 152227 79796 152293 79797
rect 152227 79732 152228 79796
rect 152292 79794 152293 79796
rect 152414 79794 152474 183499
rect 152292 79734 152474 79794
rect 152292 79732 152293 79734
rect 152227 79731 152293 79732
rect 151307 79660 151373 79661
rect 151307 79596 151308 79660
rect 151372 79596 151373 79660
rect 151307 79595 151373 79596
rect 151491 78708 151557 78709
rect 151491 78644 151492 78708
rect 151556 78644 151557 78708
rect 151491 78643 151557 78644
rect 150755 78436 150821 78437
rect 150755 78372 150756 78436
rect 150820 78372 150821 78436
rect 150755 78371 150821 78372
rect 149654 73750 149898 73810
rect 150022 78102 150450 78162
rect 151123 78164 151189 78165
rect 149467 72724 149533 72725
rect 149467 72660 149468 72724
rect 149532 72660 149533 72724
rect 149467 72659 149533 72660
rect 149470 63341 149530 72659
rect 149654 71501 149714 73750
rect 150022 72589 150082 78102
rect 151123 78100 151124 78164
rect 151188 78100 151189 78164
rect 151123 78099 151189 78100
rect 150019 72588 150085 72589
rect 150019 72524 150020 72588
rect 150084 72524 150085 72588
rect 150019 72523 150085 72524
rect 149651 71500 149717 71501
rect 149651 71436 149652 71500
rect 149716 71436 149717 71500
rect 149651 71435 149717 71436
rect 149467 63340 149533 63341
rect 149467 63276 149468 63340
rect 149532 63276 149533 63340
rect 149467 63275 149533 63276
rect 149283 42124 149349 42125
rect 149283 42060 149284 42124
rect 149348 42060 149349 42124
rect 149283 42059 149349 42060
rect 148915 32468 148981 32469
rect 148915 32404 148916 32468
rect 148980 32404 148981 32468
rect 148915 32403 148981 32404
rect 149654 18597 149714 71435
rect 150022 70410 150082 72523
rect 149838 70350 150082 70410
rect 149838 61709 149898 70350
rect 149835 61708 149901 61709
rect 149835 61644 149836 61708
rect 149900 61644 149901 61708
rect 149835 61643 149901 61644
rect 150294 43954 150914 78000
rect 151126 72861 151186 78099
rect 151123 72860 151189 72861
rect 151123 72796 151124 72860
rect 151188 72796 151189 72860
rect 151123 72795 151189 72796
rect 151126 44845 151186 72795
rect 151494 67285 151554 78643
rect 152414 78573 152474 79734
rect 152598 79525 152658 199822
rect 152779 199820 152780 199822
rect 152844 199820 152845 199884
rect 152779 199819 152845 199820
rect 153147 199884 153213 199885
rect 153147 199820 153148 199884
rect 153212 199820 153213 199884
rect 153147 199819 153213 199820
rect 153331 199884 153397 199885
rect 153331 199820 153332 199884
rect 153396 199820 153397 199884
rect 153331 199819 153397 199820
rect 153150 187710 153210 199819
rect 153334 197437 153394 199819
rect 153331 197436 153397 197437
rect 153331 197372 153332 197436
rect 153396 197372 153397 197436
rect 153331 197371 153397 197372
rect 152782 187650 153210 187710
rect 152595 79524 152661 79525
rect 152595 79460 152596 79524
rect 152660 79460 152661 79524
rect 152595 79459 152661 79460
rect 152782 79389 152842 187650
rect 153518 79797 153578 199955
rect 153883 199884 153949 199885
rect 153883 199820 153884 199884
rect 153948 199820 153949 199884
rect 153883 199819 153949 199820
rect 154803 199884 154869 199885
rect 154803 199820 154804 199884
rect 154868 199820 154869 199884
rect 154803 199819 154869 199820
rect 155539 199884 155605 199885
rect 155539 199820 155540 199884
rect 155604 199820 155605 199884
rect 155539 199819 155605 199820
rect 156091 199884 156157 199885
rect 156091 199820 156092 199884
rect 156156 199820 156157 199884
rect 156091 199819 156157 199820
rect 157379 199884 157445 199885
rect 157379 199820 157380 199884
rect 157444 199820 157445 199884
rect 157379 199819 157445 199820
rect 160507 199884 160573 199885
rect 160507 199820 160508 199884
rect 160572 199820 160573 199884
rect 160507 199819 160573 199820
rect 162347 199884 162413 199885
rect 162347 199820 162348 199884
rect 162412 199820 162413 199884
rect 162347 199819 162413 199820
rect 163451 199884 163517 199885
rect 163451 199820 163452 199884
rect 163516 199820 163517 199884
rect 163451 199819 163517 199820
rect 163635 199884 163701 199885
rect 163635 199820 163636 199884
rect 163700 199820 163701 199884
rect 163635 199819 163701 199820
rect 164371 199884 164437 199885
rect 164371 199820 164372 199884
rect 164436 199820 164437 199884
rect 164371 199819 164437 199820
rect 165107 199884 165173 199885
rect 165107 199820 165108 199884
rect 165172 199820 165173 199884
rect 165107 199819 165173 199820
rect 153886 199341 153946 199819
rect 154806 199341 154866 199819
rect 153883 199340 153949 199341
rect 153883 199276 153884 199340
rect 153948 199276 153949 199340
rect 153883 199275 153949 199276
rect 154803 199340 154869 199341
rect 154803 199276 154804 199340
rect 154868 199276 154869 199340
rect 154803 199275 154869 199276
rect 154794 192454 155414 198000
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 153699 191316 153765 191317
rect 153699 191252 153700 191316
rect 153764 191252 153765 191316
rect 153699 191251 153765 191252
rect 153515 79796 153581 79797
rect 153515 79732 153516 79796
rect 153580 79732 153581 79796
rect 153515 79731 153581 79732
rect 153702 79525 153762 191251
rect 154067 190908 154133 190909
rect 154067 190844 154068 190908
rect 154132 190844 154133 190908
rect 154067 190843 154133 190844
rect 153883 189412 153949 189413
rect 153883 189348 153884 189412
rect 153948 189348 153949 189412
rect 153883 189347 153949 189348
rect 153886 79933 153946 189347
rect 153883 79932 153949 79933
rect 153883 79868 153884 79932
rect 153948 79868 153949 79932
rect 153883 79867 153949 79868
rect 153699 79524 153765 79525
rect 153699 79460 153700 79524
rect 153764 79460 153765 79524
rect 153699 79459 153765 79460
rect 152779 79388 152845 79389
rect 152779 79324 152780 79388
rect 152844 79324 152845 79388
rect 152779 79323 152845 79324
rect 152411 78572 152477 78573
rect 152411 78508 152412 78572
rect 152476 78508 152477 78572
rect 152411 78507 152477 78508
rect 152411 78300 152477 78301
rect 152411 78236 152412 78300
rect 152476 78236 152477 78300
rect 152411 78235 152477 78236
rect 152414 71637 152474 78235
rect 152963 78164 153029 78165
rect 152963 78100 152964 78164
rect 153028 78100 153029 78164
rect 152963 78099 153029 78100
rect 152779 77892 152845 77893
rect 152779 77828 152780 77892
rect 152844 77828 152845 77892
rect 152779 77827 152845 77828
rect 152411 71636 152477 71637
rect 152411 71572 152412 71636
rect 152476 71572 152477 71636
rect 152411 71571 152477 71572
rect 151491 67284 151557 67285
rect 151491 67220 151492 67284
rect 151556 67220 151557 67284
rect 151491 67219 151557 67220
rect 151123 44844 151189 44845
rect 151123 44780 151124 44844
rect 151188 44780 151189 44844
rect 151123 44779 151189 44780
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 149651 18596 149717 18597
rect 149651 18532 149652 18596
rect 149716 18532 149717 18596
rect 149651 18531 149717 18532
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 7954 150914 43398
rect 152414 26893 152474 71571
rect 152782 57901 152842 77827
rect 152966 75717 153026 78099
rect 153702 77893 153762 79459
rect 153886 79389 153946 79867
rect 154070 79661 154130 190843
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 155355 139364 155421 139365
rect 155355 139300 155356 139364
rect 155420 139300 155421 139364
rect 155355 139299 155421 139300
rect 154803 139228 154869 139229
rect 154803 139164 154804 139228
rect 154868 139164 154869 139228
rect 154803 139163 154869 139164
rect 154806 80205 154866 139163
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 154803 80204 154869 80205
rect 154803 80140 154804 80204
rect 154868 80140 154869 80204
rect 154803 80139 154869 80140
rect 155358 79933 155418 139299
rect 155355 79932 155421 79933
rect 155355 79868 155356 79932
rect 155420 79868 155421 79932
rect 155355 79867 155421 79868
rect 155355 79796 155421 79797
rect 155355 79732 155356 79796
rect 155420 79794 155421 79796
rect 155542 79794 155602 199819
rect 156094 199341 156154 199819
rect 156827 199476 156893 199477
rect 156827 199412 156828 199476
rect 156892 199412 156893 199476
rect 156827 199411 156893 199412
rect 156091 199340 156157 199341
rect 156091 199276 156092 199340
rect 156156 199276 156157 199340
rect 156091 199275 156157 199276
rect 156643 197300 156709 197301
rect 156643 197236 156644 197300
rect 156708 197236 156709 197300
rect 156643 197235 156709 197236
rect 156275 195668 156341 195669
rect 156275 195604 156276 195668
rect 156340 195604 156341 195668
rect 156275 195603 156341 195604
rect 155723 194036 155789 194037
rect 155723 193972 155724 194036
rect 155788 193972 155789 194036
rect 155723 193971 155789 193972
rect 155726 80069 155786 193971
rect 156278 80069 156338 195603
rect 156646 80341 156706 197235
rect 156643 80340 156709 80341
rect 156643 80276 156644 80340
rect 156708 80276 156709 80340
rect 156643 80275 156709 80276
rect 155723 80068 155789 80069
rect 155723 80004 155724 80068
rect 155788 80004 155789 80068
rect 155723 80003 155789 80004
rect 156275 80068 156341 80069
rect 156275 80004 156276 80068
rect 156340 80004 156341 80068
rect 156275 80003 156341 80004
rect 155420 79734 155602 79794
rect 155420 79732 155421 79734
rect 155355 79731 155421 79732
rect 154067 79660 154133 79661
rect 154067 79596 154068 79660
rect 154132 79596 154133 79660
rect 154067 79595 154133 79596
rect 154251 79660 154317 79661
rect 154251 79596 154252 79660
rect 154316 79596 154317 79660
rect 154251 79595 154317 79596
rect 153883 79388 153949 79389
rect 153883 79324 153884 79388
rect 153948 79324 153949 79388
rect 153883 79323 153949 79324
rect 154067 78572 154133 78573
rect 154067 78508 154068 78572
rect 154132 78508 154133 78572
rect 154067 78507 154133 78508
rect 153699 77892 153765 77893
rect 153699 77828 153700 77892
rect 153764 77828 153765 77892
rect 153699 77827 153765 77828
rect 153883 76668 153949 76669
rect 153883 76604 153884 76668
rect 153948 76604 153949 76668
rect 153883 76603 153949 76604
rect 152963 75716 153029 75717
rect 152963 75652 152964 75716
rect 153028 75652 153029 75716
rect 152963 75651 153029 75652
rect 152779 57900 152845 57901
rect 152779 57836 152780 57900
rect 152844 57836 152845 57900
rect 152779 57835 152845 57836
rect 152966 40629 153026 75651
rect 153886 66197 153946 76603
rect 153883 66196 153949 66197
rect 153883 66132 153884 66196
rect 153948 66132 153949 66196
rect 153883 66131 153949 66132
rect 154070 63205 154130 78507
rect 154067 63204 154133 63205
rect 154067 63140 154068 63204
rect 154132 63140 154133 63204
rect 154067 63139 154133 63140
rect 154254 59125 154314 79595
rect 155726 79525 155786 80003
rect 156459 79932 156525 79933
rect 156459 79868 156460 79932
rect 156524 79868 156525 79932
rect 156459 79867 156525 79868
rect 155723 79524 155789 79525
rect 155723 79460 155724 79524
rect 155788 79460 155789 79524
rect 155723 79459 155789 79460
rect 154435 78572 154501 78573
rect 154435 78508 154436 78572
rect 154500 78508 154501 78572
rect 154435 78507 154501 78508
rect 155723 78572 155789 78573
rect 155723 78508 155724 78572
rect 155788 78508 155789 78572
rect 155723 78507 155789 78508
rect 154251 59124 154317 59125
rect 154251 59060 154252 59124
rect 154316 59060 154317 59124
rect 154251 59059 154317 59060
rect 154438 53549 154498 78507
rect 154435 53548 154501 53549
rect 154435 53484 154436 53548
rect 154500 53484 154501 53548
rect 154435 53483 154501 53484
rect 154794 48454 155414 78000
rect 155539 77892 155605 77893
rect 155539 77828 155540 77892
rect 155604 77828 155605 77892
rect 155539 77827 155605 77828
rect 155542 67421 155602 77827
rect 155539 67420 155605 67421
rect 155539 67356 155540 67420
rect 155604 67356 155605 67420
rect 155539 67355 155605 67356
rect 155726 63069 155786 78507
rect 156275 78164 156341 78165
rect 156275 78100 156276 78164
rect 156340 78100 156341 78164
rect 156275 78099 156341 78100
rect 156278 75930 156338 78099
rect 156462 77621 156522 79867
rect 156830 79661 156890 199411
rect 157382 199341 157442 199819
rect 157379 199340 157445 199341
rect 157379 199276 157380 199340
rect 157444 199276 157445 199340
rect 157379 199275 157445 199276
rect 158299 199340 158365 199341
rect 158299 199276 158300 199340
rect 158364 199276 158365 199340
rect 158299 199275 158365 199276
rect 157195 198932 157261 198933
rect 157195 198868 157196 198932
rect 157260 198868 157261 198932
rect 157195 198867 157261 198868
rect 157011 198796 157077 198797
rect 157011 198732 157012 198796
rect 157076 198732 157077 198796
rect 157011 198731 157077 198732
rect 157014 79797 157074 198731
rect 157198 197437 157258 198867
rect 158115 198796 158181 198797
rect 158115 198732 158116 198796
rect 158180 198732 158181 198796
rect 158115 198731 158181 198732
rect 157563 198252 157629 198253
rect 157563 198188 157564 198252
rect 157628 198188 157629 198252
rect 157563 198187 157629 198188
rect 157195 197436 157261 197437
rect 157195 197372 157196 197436
rect 157260 197372 157261 197436
rect 157195 197371 157261 197372
rect 157195 80340 157261 80341
rect 157195 80276 157196 80340
rect 157260 80276 157261 80340
rect 157195 80275 157261 80276
rect 157198 79933 157258 80275
rect 157195 79932 157261 79933
rect 157195 79868 157196 79932
rect 157260 79868 157261 79932
rect 157195 79867 157261 79868
rect 157011 79796 157077 79797
rect 157011 79732 157012 79796
rect 157076 79732 157077 79796
rect 157011 79731 157077 79732
rect 156827 79660 156893 79661
rect 156827 79596 156828 79660
rect 156892 79596 156893 79660
rect 156827 79595 156893 79596
rect 157566 79525 157626 198187
rect 157931 196756 157997 196757
rect 157931 196692 157932 196756
rect 157996 196692 157997 196756
rect 157931 196691 157997 196692
rect 157934 79933 157994 196691
rect 157931 79932 157997 79933
rect 157931 79868 157932 79932
rect 157996 79868 157997 79932
rect 157931 79867 157997 79868
rect 158118 79661 158178 198731
rect 158302 79933 158362 199275
rect 159294 196954 159914 198000
rect 160510 197709 160570 199819
rect 161243 199340 161309 199341
rect 161243 199276 161244 199340
rect 161308 199276 161309 199340
rect 161243 199275 161309 199276
rect 160507 197708 160573 197709
rect 160507 197644 160508 197708
rect 160572 197644 160573 197708
rect 160507 197643 160573 197644
rect 160875 197436 160941 197437
rect 160875 197372 160876 197436
rect 160940 197372 160941 197436
rect 160875 197371 160941 197372
rect 160507 197164 160573 197165
rect 160507 197100 160508 197164
rect 160572 197100 160573 197164
rect 160507 197099 160573 197100
rect 158851 196756 158917 196757
rect 158851 196692 158852 196756
rect 158916 196692 158917 196756
rect 158851 196691 158917 196692
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 158854 86970 158914 196691
rect 159294 196634 159914 196718
rect 159035 196620 159101 196621
rect 159035 196556 159036 196620
rect 159100 196556 159101 196620
rect 159035 196555 159101 196556
rect 158670 86910 158914 86970
rect 158299 79932 158365 79933
rect 158299 79868 158300 79932
rect 158364 79868 158365 79932
rect 158299 79867 158365 79868
rect 158670 79661 158730 86910
rect 158851 79932 158917 79933
rect 158851 79868 158852 79932
rect 158916 79868 158917 79932
rect 158851 79867 158917 79868
rect 157747 79660 157813 79661
rect 157747 79596 157748 79660
rect 157812 79596 157813 79660
rect 157747 79595 157813 79596
rect 158115 79660 158181 79661
rect 158115 79596 158116 79660
rect 158180 79596 158181 79660
rect 158115 79595 158181 79596
rect 158667 79660 158733 79661
rect 158667 79596 158668 79660
rect 158732 79596 158733 79660
rect 158667 79595 158733 79596
rect 157563 79524 157629 79525
rect 157563 79460 157564 79524
rect 157628 79460 157629 79524
rect 157563 79459 157629 79460
rect 156827 79388 156893 79389
rect 156827 79324 156828 79388
rect 156892 79324 156893 79388
rect 156827 79323 156893 79324
rect 156643 78436 156709 78437
rect 156643 78372 156644 78436
rect 156708 78372 156709 78436
rect 156643 78371 156709 78372
rect 156459 77620 156525 77621
rect 156459 77556 156460 77620
rect 156524 77556 156525 77620
rect 156459 77555 156525 77556
rect 156278 75870 156522 75930
rect 156462 74493 156522 75870
rect 156459 74492 156525 74493
rect 156459 74428 156460 74492
rect 156524 74428 156525 74492
rect 156459 74427 156525 74428
rect 155723 63068 155789 63069
rect 155723 63004 155724 63068
rect 155788 63004 155789 63068
rect 155723 63003 155789 63004
rect 156646 57629 156706 78371
rect 156830 73133 156890 79323
rect 157011 77892 157077 77893
rect 157011 77828 157012 77892
rect 157076 77828 157077 77892
rect 157011 77827 157077 77828
rect 156827 73132 156893 73133
rect 156827 73068 156828 73132
rect 156892 73068 156893 73132
rect 156827 73067 156893 73068
rect 157014 61981 157074 77827
rect 157750 77310 157810 79595
rect 158115 78708 158181 78709
rect 158115 78644 158116 78708
rect 158180 78644 158181 78708
rect 158115 78643 158181 78644
rect 158483 78708 158549 78709
rect 158483 78644 158484 78708
rect 158548 78644 158549 78708
rect 158483 78643 158549 78644
rect 157750 77250 157994 77310
rect 157011 61980 157077 61981
rect 157011 61916 157012 61980
rect 157076 61916 157077 61980
rect 157011 61915 157077 61916
rect 157934 58853 157994 77250
rect 157931 58852 157997 58853
rect 157931 58788 157932 58852
rect 157996 58788 157997 58852
rect 157931 58787 157997 58788
rect 156643 57628 156709 57629
rect 156643 57564 156644 57628
rect 156708 57564 156709 57628
rect 156643 57563 156709 57564
rect 158118 55045 158178 78643
rect 158299 77892 158365 77893
rect 158299 77828 158300 77892
rect 158364 77828 158365 77892
rect 158299 77827 158365 77828
rect 158115 55044 158181 55045
rect 158115 54980 158116 55044
rect 158180 54980 158181 55044
rect 158115 54979 158181 54980
rect 158302 50829 158362 77827
rect 158486 73677 158546 78643
rect 158483 73676 158549 73677
rect 158483 73612 158484 73676
rect 158548 73612 158549 73676
rect 158483 73611 158549 73612
rect 158299 50828 158365 50829
rect 158299 50764 158300 50828
rect 158364 50764 158365 50828
rect 158299 50763 158365 50764
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 152963 40628 153029 40629
rect 152963 40564 152964 40628
rect 153028 40564 153029 40628
rect 152963 40563 153029 40564
rect 152411 26892 152477 26893
rect 152411 26828 152412 26892
rect 152476 26828 152477 26892
rect 152411 26827 152477 26828
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 158486 11661 158546 73611
rect 158854 56405 158914 79867
rect 159038 79797 159098 196555
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 160510 190637 160570 197099
rect 160507 190636 160573 190637
rect 160507 190572 160508 190636
rect 160572 190572 160573 190636
rect 160507 190571 160573 190572
rect 160691 190500 160757 190501
rect 160691 190436 160692 190500
rect 160756 190436 160757 190500
rect 160691 190435 160757 190436
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 142000 159914 160398
rect 159219 139364 159285 139365
rect 159219 139300 159220 139364
rect 159284 139300 159285 139364
rect 159219 139299 159285 139300
rect 159955 139364 160021 139365
rect 159955 139300 159956 139364
rect 160020 139300 160021 139364
rect 159955 139299 160021 139300
rect 159222 89730 159282 139299
rect 159222 89670 159650 89730
rect 159590 80205 159650 89670
rect 159587 80204 159653 80205
rect 159587 80140 159588 80204
rect 159652 80140 159653 80204
rect 159587 80139 159653 80140
rect 159035 79796 159101 79797
rect 159035 79732 159036 79796
rect 159100 79732 159101 79796
rect 159035 79731 159101 79732
rect 159590 78709 159650 80139
rect 159958 79389 160018 139299
rect 160323 80884 160389 80885
rect 160323 80820 160324 80884
rect 160388 80820 160389 80884
rect 160323 80819 160389 80820
rect 160326 79933 160386 80819
rect 160323 79932 160389 79933
rect 160323 79868 160324 79932
rect 160388 79868 160389 79932
rect 160323 79867 160389 79868
rect 160694 79797 160754 190435
rect 160878 80341 160938 197371
rect 161059 197300 161125 197301
rect 161059 197236 161060 197300
rect 161124 197236 161125 197300
rect 161059 197235 161125 197236
rect 160875 80340 160941 80341
rect 160875 80276 160876 80340
rect 160940 80276 160941 80340
rect 160875 80275 160941 80276
rect 161062 80202 161122 197235
rect 161246 190770 161306 199275
rect 162163 197572 162229 197573
rect 162163 197508 162164 197572
rect 162228 197508 162229 197572
rect 162163 197507 162229 197508
rect 161979 196756 162045 196757
rect 161979 196692 161980 196756
rect 162044 196692 162045 196756
rect 161979 196691 162045 196692
rect 161246 190710 161490 190770
rect 161243 190636 161309 190637
rect 161243 190572 161244 190636
rect 161308 190572 161309 190636
rect 161243 190571 161309 190572
rect 161246 80477 161306 190571
rect 161430 190229 161490 190710
rect 161427 190228 161493 190229
rect 161427 190164 161428 190228
rect 161492 190164 161493 190228
rect 161427 190163 161493 190164
rect 161427 180844 161493 180845
rect 161427 180780 161428 180844
rect 161492 180780 161493 180844
rect 161427 180779 161493 180780
rect 161430 180573 161490 180779
rect 161427 180572 161493 180573
rect 161427 180508 161428 180572
rect 161492 180508 161493 180572
rect 161427 180507 161493 180508
rect 161427 171188 161493 171189
rect 161427 171124 161428 171188
rect 161492 171124 161493 171188
rect 161427 171123 161493 171124
rect 161430 170917 161490 171123
rect 161427 170916 161493 170917
rect 161427 170852 161428 170916
rect 161492 170852 161493 170916
rect 161427 170851 161493 170852
rect 161427 161532 161493 161533
rect 161427 161468 161428 161532
rect 161492 161468 161493 161532
rect 161427 161467 161493 161468
rect 161430 161261 161490 161467
rect 161427 161260 161493 161261
rect 161427 161196 161428 161260
rect 161492 161196 161493 161260
rect 161427 161195 161493 161196
rect 161427 151876 161493 151877
rect 161427 151812 161428 151876
rect 161492 151812 161493 151876
rect 161427 151811 161493 151812
rect 161430 151605 161490 151811
rect 161427 151604 161493 151605
rect 161427 151540 161428 151604
rect 161492 151540 161493 151604
rect 161427 151539 161493 151540
rect 161611 142356 161677 142357
rect 161611 142292 161612 142356
rect 161676 142292 161677 142356
rect 161611 142291 161677 142292
rect 161243 80476 161309 80477
rect 161243 80412 161244 80476
rect 161308 80412 161309 80476
rect 161243 80411 161309 80412
rect 160878 80142 161122 80202
rect 160691 79796 160757 79797
rect 160691 79732 160692 79796
rect 160756 79732 160757 79796
rect 160691 79731 160757 79732
rect 160878 79661 160938 80142
rect 161427 79932 161493 79933
rect 161427 79868 161428 79932
rect 161492 79868 161493 79932
rect 161427 79867 161493 79868
rect 160875 79660 160941 79661
rect 160875 79596 160876 79660
rect 160940 79596 160941 79660
rect 160875 79595 160941 79596
rect 159955 79388 160021 79389
rect 159955 79324 159956 79388
rect 160020 79324 160021 79388
rect 159955 79323 160021 79324
rect 160691 79116 160757 79117
rect 160691 79052 160692 79116
rect 160756 79052 160757 79116
rect 160691 79051 160757 79052
rect 159587 78708 159653 78709
rect 159587 78644 159588 78708
rect 159652 78644 159653 78708
rect 159587 78643 159653 78644
rect 159035 78436 159101 78437
rect 159035 78372 159036 78436
rect 159100 78372 159101 78436
rect 159035 78371 159101 78372
rect 158851 56404 158917 56405
rect 158851 56340 158852 56404
rect 158916 56340 158917 56404
rect 158851 56339 158917 56340
rect 159038 49333 159098 78371
rect 159294 52954 159914 78000
rect 160694 66061 160754 79051
rect 160875 77348 160941 77349
rect 160875 77284 160876 77348
rect 160940 77284 160941 77348
rect 160875 77283 160941 77284
rect 161059 77348 161125 77349
rect 161059 77284 161060 77348
rect 161124 77284 161125 77348
rect 161059 77283 161125 77284
rect 160691 66060 160757 66061
rect 160691 65996 160692 66060
rect 160756 65996 160757 66060
rect 160691 65995 160757 65996
rect 160878 57493 160938 77283
rect 160875 57492 160941 57493
rect 160875 57428 160876 57492
rect 160940 57428 160941 57492
rect 160875 57427 160941 57428
rect 161062 54909 161122 77283
rect 161430 73170 161490 79867
rect 161614 79525 161674 142291
rect 161982 80069 162042 196691
rect 161979 80068 162045 80069
rect 161979 80004 161980 80068
rect 162044 80004 162045 80068
rect 161979 80003 162045 80004
rect 162166 79933 162226 197507
rect 162163 79932 162229 79933
rect 162163 79868 162164 79932
rect 162228 79868 162229 79932
rect 162163 79867 162229 79868
rect 162163 79660 162229 79661
rect 162163 79596 162164 79660
rect 162228 79596 162229 79660
rect 162163 79595 162229 79596
rect 161611 79524 161677 79525
rect 161611 79460 161612 79524
rect 161676 79460 161677 79524
rect 161611 79459 161677 79460
rect 161246 73110 161490 73170
rect 161059 54908 161125 54909
rect 161059 54844 161060 54908
rect 161124 54844 161125 54908
rect 161059 54843 161125 54844
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159035 49332 159101 49333
rect 159035 49268 159036 49332
rect 159100 49268 159101 49332
rect 159035 49267 159101 49268
rect 159294 16954 159914 52398
rect 161246 48109 161306 73110
rect 162166 66741 162226 79595
rect 162350 79525 162410 199819
rect 163083 197436 163149 197437
rect 163083 197372 163084 197436
rect 163148 197372 163149 197436
rect 163083 197371 163149 197372
rect 163086 79661 163146 197371
rect 163267 197300 163333 197301
rect 163267 197236 163268 197300
rect 163332 197236 163333 197300
rect 163267 197235 163333 197236
rect 163083 79660 163149 79661
rect 163083 79596 163084 79660
rect 163148 79596 163149 79660
rect 163083 79595 163149 79596
rect 163270 79525 163330 197235
rect 163454 191181 163514 199819
rect 163451 191180 163517 191181
rect 163451 191116 163452 191180
rect 163516 191116 163517 191180
rect 163451 191115 163517 191116
rect 163451 79932 163517 79933
rect 163451 79868 163452 79932
rect 163516 79868 163517 79932
rect 163451 79867 163517 79868
rect 162347 79524 162413 79525
rect 162347 79460 162348 79524
rect 162412 79460 162413 79524
rect 162347 79459 162413 79460
rect 163267 79524 163333 79525
rect 163267 79460 163268 79524
rect 163332 79460 163333 79524
rect 163267 79459 163333 79460
rect 162531 79116 162597 79117
rect 162531 79052 162532 79116
rect 162596 79052 162597 79116
rect 162531 79051 162597 79052
rect 162534 77210 162594 79051
rect 162350 77150 162594 77210
rect 162163 66740 162229 66741
rect 162163 66676 162164 66740
rect 162228 66676 162229 66740
rect 162163 66675 162229 66676
rect 162350 58717 162410 77150
rect 162531 76532 162597 76533
rect 162531 76468 162532 76532
rect 162596 76468 162597 76532
rect 163454 76530 163514 79867
rect 163638 79661 163698 199819
rect 164374 191181 164434 199819
rect 165110 199341 165170 199819
rect 165107 199340 165173 199341
rect 165107 199276 165108 199340
rect 165172 199276 165173 199340
rect 165107 199275 165173 199276
rect 164555 197572 164621 197573
rect 164555 197508 164556 197572
rect 164620 197508 164621 197572
rect 164555 197507 164621 197508
rect 164371 191180 164437 191181
rect 164371 191116 164372 191180
rect 164436 191116 164437 191180
rect 164371 191115 164437 191116
rect 164003 189412 164069 189413
rect 164003 189348 164004 189412
rect 164068 189348 164069 189412
rect 164003 189347 164069 189348
rect 163635 79660 163701 79661
rect 163635 79596 163636 79660
rect 163700 79596 163701 79660
rect 163635 79595 163701 79596
rect 164006 79253 164066 189347
rect 164187 80612 164253 80613
rect 164187 80548 164188 80612
rect 164252 80548 164253 80612
rect 164187 80547 164253 80548
rect 164190 79661 164250 80547
rect 164187 79660 164253 79661
rect 164187 79596 164188 79660
rect 164252 79596 164253 79660
rect 164187 79595 164253 79596
rect 164558 79525 164618 197507
rect 164923 197436 164989 197437
rect 164923 197372 164924 197436
rect 164988 197372 164989 197436
rect 164923 197371 164989 197372
rect 164739 191180 164805 191181
rect 164739 191116 164740 191180
rect 164804 191116 164805 191180
rect 164739 191115 164805 191116
rect 164742 79797 164802 191115
rect 164739 79796 164805 79797
rect 164739 79732 164740 79796
rect 164804 79732 164805 79796
rect 164739 79731 164805 79732
rect 164555 79524 164621 79525
rect 164555 79460 164556 79524
rect 164620 79460 164621 79524
rect 164555 79459 164621 79460
rect 164926 79253 164986 197371
rect 165294 197301 165354 199955
rect 166579 199884 166645 199885
rect 166579 199882 166580 199884
rect 166030 199822 166580 199882
rect 166030 198933 166090 199822
rect 166579 199820 166580 199822
rect 166644 199820 166645 199884
rect 166579 199819 166645 199820
rect 167131 199884 167197 199885
rect 167131 199820 167132 199884
rect 167196 199820 167197 199884
rect 167545 199884 167611 199885
rect 167545 199882 167546 199884
rect 167131 199819 167197 199820
rect 167502 199820 167546 199882
rect 167610 199820 167611 199884
rect 167502 199819 167611 199820
rect 167867 199884 167933 199885
rect 167867 199820 167868 199884
rect 167932 199820 167933 199884
rect 167867 199819 167933 199820
rect 166395 199068 166461 199069
rect 166395 199004 166396 199068
rect 166460 199004 166461 199068
rect 166395 199003 166461 199004
rect 166027 198932 166093 198933
rect 166027 198868 166028 198932
rect 166092 198868 166093 198932
rect 166027 198867 166093 198868
rect 166211 198932 166277 198933
rect 166211 198868 166212 198932
rect 166276 198868 166277 198932
rect 166211 198867 166277 198868
rect 165107 197300 165173 197301
rect 165107 197236 165108 197300
rect 165172 197236 165173 197300
rect 165107 197235 165173 197236
rect 165291 197300 165357 197301
rect 165291 197236 165292 197300
rect 165356 197236 165357 197300
rect 165291 197235 165357 197236
rect 165659 197300 165725 197301
rect 165659 197236 165660 197300
rect 165724 197236 165725 197300
rect 165659 197235 165725 197236
rect 165110 79797 165170 197235
rect 165662 89730 165722 197235
rect 165662 89670 165906 89730
rect 165475 80068 165541 80069
rect 165475 80004 165476 80068
rect 165540 80004 165541 80068
rect 165475 80003 165541 80004
rect 165291 79932 165357 79933
rect 165291 79868 165292 79932
rect 165356 79868 165357 79932
rect 165291 79867 165357 79868
rect 165107 79796 165173 79797
rect 165107 79732 165108 79796
rect 165172 79732 165173 79796
rect 165107 79731 165173 79732
rect 164003 79252 164069 79253
rect 164003 79188 164004 79252
rect 164068 79188 164069 79252
rect 164003 79187 164069 79188
rect 164923 79252 164989 79253
rect 164923 79188 164924 79252
rect 164988 79188 164989 79252
rect 164923 79187 164989 79188
rect 163454 76470 163698 76530
rect 162531 76467 162597 76468
rect 162347 58716 162413 58717
rect 162347 58652 162348 58716
rect 162412 58652 162413 58716
rect 162347 58651 162413 58652
rect 162534 53685 162594 76467
rect 163267 76124 163333 76125
rect 163267 76060 163268 76124
rect 163332 76060 163333 76124
rect 163267 76059 163333 76060
rect 162715 75988 162781 75989
rect 162715 75924 162716 75988
rect 162780 75924 162781 75988
rect 162715 75923 162781 75924
rect 162531 53684 162597 53685
rect 162531 53620 162532 53684
rect 162596 53620 162597 53684
rect 162531 53619 162597 53620
rect 162718 49469 162778 75923
rect 163270 56269 163330 76059
rect 163451 75988 163517 75989
rect 163451 75924 163452 75988
rect 163516 75924 163517 75988
rect 163451 75923 163517 75924
rect 163267 56268 163333 56269
rect 163267 56204 163268 56268
rect 163332 56204 163333 56268
rect 163267 56203 163333 56204
rect 163454 55181 163514 75923
rect 163451 55180 163517 55181
rect 163451 55116 163452 55180
rect 163516 55116 163517 55180
rect 163451 55115 163517 55116
rect 163638 52325 163698 76470
rect 163794 57454 164414 78000
rect 165294 77890 165354 79867
rect 164926 77830 165354 77890
rect 164926 61845 164986 77830
rect 165107 77620 165173 77621
rect 165107 77556 165108 77620
rect 165172 77556 165173 77620
rect 165107 77555 165173 77556
rect 164923 61844 164989 61845
rect 164923 61780 164924 61844
rect 164988 61780 164989 61844
rect 164923 61779 164989 61780
rect 165110 60621 165170 77555
rect 165478 76530 165538 80003
rect 165846 79661 165906 89670
rect 166027 79796 166093 79797
rect 166027 79732 166028 79796
rect 166092 79732 166093 79796
rect 166027 79731 166093 79732
rect 165843 79660 165909 79661
rect 165843 79596 165844 79660
rect 165908 79596 165909 79660
rect 165843 79595 165909 79596
rect 165294 76470 165538 76530
rect 165107 60620 165173 60621
rect 165107 60556 165108 60620
rect 165172 60556 165173 60620
rect 165107 60555 165173 60556
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 165294 57357 165354 76470
rect 165475 76124 165541 76125
rect 165475 76060 165476 76124
rect 165540 76060 165541 76124
rect 165475 76059 165541 76060
rect 165291 57356 165357 57357
rect 165291 57292 165292 57356
rect 165356 57292 165357 57356
rect 165291 57291 165357 57292
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163635 52324 163701 52325
rect 163635 52260 163636 52324
rect 163700 52260 163701 52324
rect 163635 52259 163701 52260
rect 162715 49468 162781 49469
rect 162715 49404 162716 49468
rect 162780 49404 162781 49468
rect 162715 49403 162781 49404
rect 161243 48108 161309 48109
rect 161243 48044 161244 48108
rect 161308 48044 161309 48108
rect 161243 48043 161309 48044
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 158483 11660 158549 11661
rect 158483 11596 158484 11660
rect 158548 11596 158549 11660
rect 158483 11595 158549 11596
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 21454 164414 56898
rect 165478 50965 165538 76059
rect 166030 71790 166090 79731
rect 166214 79253 166274 198867
rect 166398 80069 166458 199003
rect 166579 198116 166645 198117
rect 166579 198052 166580 198116
rect 166644 198052 166645 198116
rect 166579 198051 166645 198052
rect 166395 80068 166461 80069
rect 166395 80004 166396 80068
rect 166460 80004 166461 80068
rect 166395 80003 166461 80004
rect 166211 79252 166277 79253
rect 166211 79188 166212 79252
rect 166276 79188 166277 79252
rect 166211 79187 166277 79188
rect 166398 78029 166458 80003
rect 166582 79933 166642 198051
rect 167134 193221 167194 199819
rect 167315 197300 167381 197301
rect 167315 197236 167316 197300
rect 167380 197236 167381 197300
rect 167315 197235 167381 197236
rect 167131 193220 167197 193221
rect 167131 193156 167132 193220
rect 167196 193156 167197 193220
rect 167131 193155 167197 193156
rect 167318 80205 167378 197235
rect 167315 80204 167381 80205
rect 167315 80140 167316 80204
rect 167380 80140 167381 80204
rect 167315 80139 167381 80140
rect 166579 79932 166645 79933
rect 166579 79868 166580 79932
rect 166644 79868 166645 79932
rect 166579 79867 166645 79868
rect 166947 79932 167013 79933
rect 166947 79868 166948 79932
rect 167012 79868 167013 79932
rect 167502 79930 167562 199819
rect 167870 198933 167930 199819
rect 167867 198932 167933 198933
rect 167867 198868 167868 198932
rect 167932 198868 167933 198932
rect 167867 198867 167933 198868
rect 167683 197572 167749 197573
rect 167683 197508 167684 197572
rect 167748 197508 167749 197572
rect 167683 197507 167749 197508
rect 166947 79867 167013 79868
rect 167318 79870 167562 79930
rect 166763 79524 166829 79525
rect 166763 79460 166764 79524
rect 166828 79460 166829 79524
rect 166763 79459 166829 79460
rect 166395 78028 166461 78029
rect 166395 77964 166396 78028
rect 166460 77964 166461 78028
rect 166395 77963 166461 77964
rect 166395 75988 166461 75989
rect 166395 75924 166396 75988
rect 166460 75924 166461 75988
rect 166395 75923 166461 75924
rect 166579 75988 166645 75989
rect 166579 75924 166580 75988
rect 166644 75924 166645 75988
rect 166579 75923 166645 75924
rect 166030 71730 166274 71790
rect 166214 63477 166274 71730
rect 166211 63476 166277 63477
rect 166211 63412 166212 63476
rect 166276 63412 166277 63476
rect 166211 63411 166277 63412
rect 166398 53821 166458 75923
rect 166395 53820 166461 53821
rect 166395 53756 166396 53820
rect 166460 53756 166461 53820
rect 166395 53755 166461 53756
rect 165475 50964 165541 50965
rect 165475 50900 165476 50964
rect 165540 50900 165541 50964
rect 165475 50899 165541 50900
rect 166582 49605 166642 75923
rect 166579 49604 166645 49605
rect 166579 49540 166580 49604
rect 166644 49540 166645 49604
rect 166579 49539 166645 49540
rect 166766 44165 166826 79459
rect 166950 79117 167010 79867
rect 167318 79525 167378 79870
rect 167499 79796 167565 79797
rect 167499 79732 167500 79796
rect 167564 79732 167565 79796
rect 167499 79731 167565 79732
rect 167315 79524 167381 79525
rect 167315 79460 167316 79524
rect 167380 79460 167381 79524
rect 167315 79459 167381 79460
rect 166947 79116 167013 79117
rect 166947 79052 166948 79116
rect 167012 79052 167013 79116
rect 166947 79051 167013 79052
rect 167502 59261 167562 79731
rect 167686 79525 167746 197507
rect 168051 197436 168117 197437
rect 168051 197372 168052 197436
rect 168116 197372 168117 197436
rect 168051 197371 168117 197372
rect 168054 84210 168114 197371
rect 168790 196621 168850 199955
rect 168971 199884 169037 199885
rect 168971 199820 168972 199884
rect 169036 199820 169037 199884
rect 168971 199819 169037 199820
rect 168787 196620 168853 196621
rect 168787 196556 168788 196620
rect 168852 196556 168853 196620
rect 168787 196555 168853 196556
rect 167870 84150 168114 84210
rect 167870 79661 167930 84150
rect 168603 80068 168669 80069
rect 168603 80004 168604 80068
rect 168668 80004 168669 80068
rect 168603 80003 168669 80004
rect 168051 79932 168117 79933
rect 168051 79868 168052 79932
rect 168116 79868 168117 79932
rect 168051 79867 168117 79868
rect 168235 79932 168301 79933
rect 168235 79868 168236 79932
rect 168300 79868 168301 79932
rect 168235 79867 168301 79868
rect 167867 79660 167933 79661
rect 167867 79596 167868 79660
rect 167932 79596 167933 79660
rect 167867 79595 167933 79596
rect 167683 79524 167749 79525
rect 167683 79460 167684 79524
rect 167748 79460 167749 79524
rect 167683 79459 167749 79460
rect 167867 79116 167933 79117
rect 167867 79052 167868 79116
rect 167932 79052 167933 79116
rect 167867 79051 167933 79052
rect 167683 75988 167749 75989
rect 167683 75924 167684 75988
rect 167748 75924 167749 75988
rect 167683 75923 167749 75924
rect 167499 59260 167565 59261
rect 167499 59196 167500 59260
rect 167564 59196 167565 59260
rect 167499 59195 167565 59196
rect 167686 56541 167746 75923
rect 167683 56540 167749 56541
rect 167683 56476 167684 56540
rect 167748 56476 167749 56540
rect 167683 56475 167749 56476
rect 167870 52461 167930 79051
rect 167867 52460 167933 52461
rect 167867 52396 167868 52460
rect 167932 52396 167933 52460
rect 167867 52395 167933 52396
rect 168054 46885 168114 79867
rect 168238 78709 168298 79867
rect 168235 78708 168301 78709
rect 168235 78644 168236 78708
rect 168300 78644 168301 78708
rect 168235 78643 168301 78644
rect 168606 78301 168666 80003
rect 168974 79117 169034 199819
rect 170262 199341 170322 200227
rect 174675 200020 174741 200021
rect 174675 199956 174676 200020
rect 174740 199956 174741 200020
rect 174675 199955 174741 199956
rect 170811 199884 170877 199885
rect 170811 199820 170812 199884
rect 170876 199882 170877 199884
rect 171363 199884 171429 199885
rect 170876 199822 171058 199882
rect 170876 199820 170877 199822
rect 170811 199819 170877 199820
rect 170259 199340 170325 199341
rect 170259 199276 170260 199340
rect 170324 199276 170325 199340
rect 170259 199275 170325 199276
rect 170443 199340 170509 199341
rect 170443 199276 170444 199340
rect 170508 199276 170509 199340
rect 170443 199275 170509 199276
rect 170811 199340 170877 199341
rect 170811 199276 170812 199340
rect 170876 199276 170877 199340
rect 170811 199275 170877 199276
rect 169891 198252 169957 198253
rect 169891 198188 169892 198252
rect 169956 198188 169957 198252
rect 169891 198187 169957 198188
rect 169155 197980 169221 197981
rect 169155 197916 169156 197980
rect 169220 197916 169221 197980
rect 169155 197915 169221 197916
rect 169158 79661 169218 197915
rect 169523 197436 169589 197437
rect 169523 197372 169524 197436
rect 169588 197372 169589 197436
rect 169523 197371 169589 197372
rect 169339 197300 169405 197301
rect 169339 197236 169340 197300
rect 169404 197236 169405 197300
rect 169339 197235 169405 197236
rect 169342 79797 169402 197235
rect 169339 79796 169405 79797
rect 169339 79732 169340 79796
rect 169404 79732 169405 79796
rect 169339 79731 169405 79732
rect 169155 79660 169221 79661
rect 169155 79596 169156 79660
rect 169220 79596 169221 79660
rect 169155 79595 169221 79596
rect 169526 79525 169586 197371
rect 169894 79797 169954 198187
rect 170075 197436 170141 197437
rect 170075 197372 170076 197436
rect 170140 197372 170141 197436
rect 170075 197371 170141 197372
rect 169707 79796 169773 79797
rect 169707 79732 169708 79796
rect 169772 79732 169773 79796
rect 169707 79731 169773 79732
rect 169891 79796 169957 79797
rect 169891 79732 169892 79796
rect 169956 79732 169957 79796
rect 169891 79731 169957 79732
rect 169523 79524 169589 79525
rect 169523 79460 169524 79524
rect 169588 79460 169589 79524
rect 169523 79459 169589 79460
rect 168971 79116 169037 79117
rect 168971 79052 168972 79116
rect 169036 79052 169037 79116
rect 168971 79051 169037 79052
rect 168603 78300 168669 78301
rect 168603 78236 168604 78300
rect 168668 78236 168669 78300
rect 168603 78235 168669 78236
rect 168294 61954 168914 78000
rect 169339 76940 169405 76941
rect 169339 76876 169340 76940
rect 169404 76876 169405 76940
rect 169339 76875 169405 76876
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 168051 46884 168117 46885
rect 168051 46820 168052 46884
rect 168116 46820 168117 46884
rect 168051 46819 168117 46820
rect 166763 44164 166829 44165
rect 166763 44100 166764 44164
rect 166828 44100 166829 44164
rect 166763 44099 166829 44100
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 61398
rect 169342 48245 169402 76875
rect 169710 75930 169770 79731
rect 170078 79661 170138 197371
rect 170446 197301 170506 199275
rect 170443 197300 170509 197301
rect 170443 197236 170444 197300
rect 170508 197236 170509 197300
rect 170443 197235 170509 197236
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 170443 80748 170509 80749
rect 170443 80684 170444 80748
rect 170508 80684 170509 80748
rect 170443 80683 170509 80684
rect 170259 80204 170325 80205
rect 170259 80140 170260 80204
rect 170324 80140 170325 80204
rect 170259 80139 170325 80140
rect 170075 79660 170141 79661
rect 170075 79596 170076 79660
rect 170140 79596 170141 79660
rect 170075 79595 170141 79596
rect 170262 76669 170322 80139
rect 170446 79389 170506 80683
rect 170627 80340 170693 80341
rect 170627 80276 170628 80340
rect 170692 80276 170693 80340
rect 170627 80275 170693 80276
rect 170630 79525 170690 80275
rect 170627 79524 170693 79525
rect 170627 79460 170628 79524
rect 170692 79460 170693 79524
rect 170627 79459 170693 79460
rect 170443 79388 170509 79389
rect 170443 79324 170444 79388
rect 170508 79324 170509 79388
rect 170443 79323 170509 79324
rect 170814 79117 170874 199275
rect 170998 79933 171058 199822
rect 171363 199820 171364 199884
rect 171428 199820 171429 199884
rect 171363 199819 171429 199820
rect 171547 199884 171613 199885
rect 171547 199820 171548 199884
rect 171612 199820 171613 199884
rect 171547 199819 171613 199820
rect 172467 199884 172533 199885
rect 172467 199820 172468 199884
rect 172532 199820 172533 199884
rect 172467 199819 172533 199820
rect 172651 199884 172717 199885
rect 172651 199820 172652 199884
rect 172716 199820 172717 199884
rect 172651 199819 172717 199820
rect 174491 199884 174557 199885
rect 174491 199820 174492 199884
rect 174556 199820 174557 199884
rect 174491 199819 174557 199820
rect 171366 199341 171426 199819
rect 171363 199340 171429 199341
rect 171363 199276 171364 199340
rect 171428 199276 171429 199340
rect 171363 199275 171429 199276
rect 171363 197436 171429 197437
rect 171363 197372 171364 197436
rect 171428 197372 171429 197436
rect 171363 197371 171429 197372
rect 170995 79932 171061 79933
rect 170995 79868 170996 79932
rect 171060 79868 171061 79932
rect 170995 79867 171061 79868
rect 170811 79116 170877 79117
rect 170811 79052 170812 79116
rect 170876 79052 170877 79116
rect 170811 79051 170877 79052
rect 170259 76668 170325 76669
rect 170259 76604 170260 76668
rect 170324 76604 170325 76668
rect 170259 76603 170325 76604
rect 170814 76533 170874 79051
rect 170998 78981 171058 79867
rect 171179 79796 171245 79797
rect 171179 79732 171180 79796
rect 171244 79732 171245 79796
rect 171179 79731 171245 79732
rect 170995 78980 171061 78981
rect 170995 78916 170996 78980
rect 171060 78916 171061 78980
rect 170995 78915 171061 78916
rect 170995 77620 171061 77621
rect 170995 77556 170996 77620
rect 171060 77556 171061 77620
rect 170995 77555 171061 77556
rect 170811 76532 170877 76533
rect 170811 76468 170812 76532
rect 170876 76468 170877 76532
rect 170811 76467 170877 76468
rect 169526 75870 169770 75930
rect 169339 48244 169405 48245
rect 169339 48180 169340 48244
rect 169404 48180 169405 48244
rect 169339 48179 169405 48180
rect 169526 44029 169586 75870
rect 170998 75173 171058 77555
rect 171182 75309 171242 79731
rect 171366 79661 171426 197371
rect 171550 79933 171610 199819
rect 171731 199340 171797 199341
rect 171731 199276 171732 199340
rect 171796 199276 171797 199340
rect 171731 199275 171797 199276
rect 171734 79933 171794 199275
rect 172470 198797 172530 199819
rect 172467 198796 172533 198797
rect 172467 198732 172468 198796
rect 172532 198732 172533 198796
rect 172467 198731 172533 198732
rect 171915 197436 171981 197437
rect 171915 197372 171916 197436
rect 171980 197372 171981 197436
rect 171915 197371 171981 197372
rect 171547 79932 171613 79933
rect 171547 79868 171548 79932
rect 171612 79868 171613 79932
rect 171547 79867 171613 79868
rect 171731 79932 171797 79933
rect 171731 79868 171732 79932
rect 171796 79868 171797 79932
rect 171731 79867 171797 79868
rect 171363 79660 171429 79661
rect 171363 79596 171364 79660
rect 171428 79596 171429 79660
rect 171363 79595 171429 79596
rect 171550 78301 171610 79867
rect 171547 78300 171613 78301
rect 171547 78236 171548 78300
rect 171612 78236 171613 78300
rect 171547 78235 171613 78236
rect 171734 77621 171794 79867
rect 171918 79253 171978 197371
rect 172099 79796 172165 79797
rect 172099 79732 172100 79796
rect 172164 79794 172165 79796
rect 172164 79734 172346 79794
rect 172164 79732 172165 79734
rect 172099 79731 172165 79732
rect 171915 79252 171981 79253
rect 171915 79188 171916 79252
rect 171980 79188 171981 79252
rect 171915 79187 171981 79188
rect 172099 78980 172165 78981
rect 172099 78916 172100 78980
rect 172164 78916 172165 78980
rect 172099 78915 172165 78916
rect 171915 78572 171981 78573
rect 171915 78508 171916 78572
rect 171980 78508 171981 78572
rect 171915 78507 171981 78508
rect 171731 77620 171797 77621
rect 171731 77556 171732 77620
rect 171796 77556 171797 77620
rect 171731 77555 171797 77556
rect 171179 75308 171245 75309
rect 171179 75244 171180 75308
rect 171244 75244 171245 75308
rect 171179 75243 171245 75244
rect 170995 75172 171061 75173
rect 170995 75108 170996 75172
rect 171060 75108 171061 75172
rect 170995 75107 171061 75108
rect 169523 44028 169589 44029
rect 169523 43964 169524 44028
rect 169588 43964 169589 44028
rect 169523 43963 169589 43964
rect 170998 36549 171058 75107
rect 171918 65789 171978 78507
rect 171915 65788 171981 65789
rect 171915 65724 171916 65788
rect 171980 65724 171981 65788
rect 171915 65723 171981 65724
rect 172102 64701 172162 78915
rect 172099 64700 172165 64701
rect 172099 64636 172100 64700
rect 172164 64636 172165 64700
rect 172099 64635 172165 64636
rect 172286 55997 172346 79734
rect 172654 79525 172714 199819
rect 174494 199477 174554 199819
rect 174678 199477 174738 199955
rect 175043 199884 175109 199885
rect 175043 199820 175044 199884
rect 175108 199820 175109 199884
rect 175043 199819 175109 199820
rect 175595 199884 175661 199885
rect 175595 199820 175596 199884
rect 175660 199820 175661 199884
rect 175595 199819 175661 199820
rect 176331 199884 176397 199885
rect 176331 199820 176332 199884
rect 176396 199820 176397 199884
rect 176331 199819 176397 199820
rect 174491 199476 174557 199477
rect 174491 199412 174492 199476
rect 174556 199412 174557 199476
rect 174491 199411 174557 199412
rect 174675 199476 174741 199477
rect 174675 199412 174676 199476
rect 174740 199412 174741 199476
rect 174675 199411 174741 199412
rect 174123 197980 174189 197981
rect 174123 197916 174124 197980
rect 174188 197916 174189 197980
rect 174123 197915 174189 197916
rect 174491 197980 174557 197981
rect 174491 197916 174492 197980
rect 174556 197916 174557 197980
rect 174491 197915 174557 197916
rect 172835 197436 172901 197437
rect 172835 197372 172836 197436
rect 172900 197372 172901 197436
rect 172835 197371 172901 197372
rect 172838 80205 172898 197371
rect 173019 197300 173085 197301
rect 173019 197236 173020 197300
rect 173084 197236 173085 197300
rect 173019 197235 173085 197236
rect 173387 197300 173453 197301
rect 173387 197236 173388 197300
rect 173452 197236 173453 197300
rect 173387 197235 173453 197236
rect 172835 80204 172901 80205
rect 172835 80140 172836 80204
rect 172900 80140 172901 80204
rect 172835 80139 172901 80140
rect 173022 79933 173082 197235
rect 173203 81156 173269 81157
rect 173203 81092 173204 81156
rect 173268 81092 173269 81156
rect 173203 81091 173269 81092
rect 173019 79932 173085 79933
rect 173019 79868 173020 79932
rect 173084 79868 173085 79932
rect 173019 79867 173085 79868
rect 173019 79796 173085 79797
rect 173019 79732 173020 79796
rect 173084 79732 173085 79796
rect 173019 79731 173085 79732
rect 172651 79524 172717 79525
rect 172651 79460 172652 79524
rect 172716 79460 172717 79524
rect 172651 79459 172717 79460
rect 173022 78437 173082 79731
rect 173206 79117 173266 81091
rect 173390 79661 173450 197235
rect 174126 79797 174186 197915
rect 174307 197436 174373 197437
rect 174307 197372 174308 197436
rect 174372 197372 174373 197436
rect 174307 197371 174373 197372
rect 173571 79796 173637 79797
rect 173571 79732 173572 79796
rect 173636 79794 173637 79796
rect 174123 79796 174189 79797
rect 173636 79734 173818 79794
rect 173636 79732 173637 79734
rect 173571 79731 173637 79732
rect 173387 79660 173453 79661
rect 173387 79596 173388 79660
rect 173452 79596 173453 79660
rect 173387 79595 173453 79596
rect 173203 79116 173269 79117
rect 173203 79052 173204 79116
rect 173268 79052 173269 79116
rect 173203 79051 173269 79052
rect 173390 78573 173450 79595
rect 173387 78572 173453 78573
rect 173387 78508 173388 78572
rect 173452 78508 173453 78572
rect 173387 78507 173453 78508
rect 173019 78436 173085 78437
rect 173019 78372 173020 78436
rect 173084 78372 173085 78436
rect 173019 78371 173085 78372
rect 172794 66454 173414 78000
rect 173571 75988 173637 75989
rect 173571 75924 173572 75988
rect 173636 75924 173637 75988
rect 173571 75923 173637 75924
rect 173574 71637 173634 75923
rect 173571 71636 173637 71637
rect 173571 71572 173572 71636
rect 173636 71572 173637 71636
rect 173571 71571 173637 71572
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172283 55996 172349 55997
rect 172283 55932 172284 55996
rect 172348 55932 172349 55996
rect 172283 55931 172349 55932
rect 170995 36548 171061 36549
rect 170995 36484 170996 36548
rect 171060 36484 171061 36548
rect 170995 36483 171061 36484
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 65898
rect 173758 65517 173818 79734
rect 174123 79732 174124 79796
rect 174188 79732 174189 79796
rect 174123 79731 174189 79732
rect 174310 79661 174370 197371
rect 174494 79794 174554 197915
rect 174859 197572 174925 197573
rect 174859 197508 174860 197572
rect 174924 197508 174925 197572
rect 174859 197507 174925 197508
rect 174862 79933 174922 197507
rect 175046 197301 175106 199819
rect 175598 199477 175658 199819
rect 175595 199476 175661 199477
rect 175595 199412 175596 199476
rect 175660 199412 175661 199476
rect 175595 199411 175661 199412
rect 175963 199068 176029 199069
rect 175963 199004 175964 199068
rect 176028 199004 176029 199068
rect 175963 199003 176029 199004
rect 175595 198524 175661 198525
rect 175595 198460 175596 198524
rect 175660 198460 175661 198524
rect 175595 198459 175661 198460
rect 175411 197436 175477 197437
rect 175411 197372 175412 197436
rect 175476 197372 175477 197436
rect 175411 197371 175477 197372
rect 175043 197300 175109 197301
rect 175043 197236 175044 197300
rect 175108 197236 175109 197300
rect 175043 197235 175109 197236
rect 175227 81020 175293 81021
rect 175227 80956 175228 81020
rect 175292 80956 175293 81020
rect 175227 80955 175293 80956
rect 174859 79932 174925 79933
rect 174859 79868 174860 79932
rect 174924 79868 174925 79932
rect 174859 79867 174925 79868
rect 175043 79932 175109 79933
rect 175043 79868 175044 79932
rect 175108 79868 175109 79932
rect 175043 79867 175109 79868
rect 174675 79796 174741 79797
rect 174675 79794 174676 79796
rect 174494 79734 174676 79794
rect 174307 79660 174373 79661
rect 174307 79596 174308 79660
rect 174372 79596 174373 79660
rect 174307 79595 174373 79596
rect 174494 77621 174554 79734
rect 174675 79732 174676 79734
rect 174740 79732 174741 79796
rect 174675 79731 174741 79732
rect 174862 78573 174922 79867
rect 174859 78572 174925 78573
rect 174859 78508 174860 78572
rect 174924 78508 174925 78572
rect 174859 78507 174925 78508
rect 174491 77620 174557 77621
rect 174491 77556 174492 77620
rect 174556 77556 174557 77620
rect 174491 77555 174557 77556
rect 174859 76940 174925 76941
rect 174859 76876 174860 76940
rect 174924 76876 174925 76940
rect 174859 76875 174925 76876
rect 174675 75580 174741 75581
rect 174675 75516 174676 75580
rect 174740 75516 174741 75580
rect 174675 75515 174741 75516
rect 173755 65516 173821 65517
rect 173755 65452 173756 65516
rect 173820 65452 173821 65516
rect 173755 65451 173821 65452
rect 174678 64837 174738 75515
rect 174675 64836 174741 64837
rect 174675 64772 174676 64836
rect 174740 64772 174741 64836
rect 174675 64771 174741 64772
rect 174862 62933 174922 76875
rect 174859 62932 174925 62933
rect 174859 62868 174860 62932
rect 174924 62868 174925 62932
rect 174859 62867 174925 62868
rect 175046 57221 175106 79867
rect 175230 79253 175290 80955
rect 175414 79525 175474 197371
rect 175598 80205 175658 198459
rect 175779 197300 175845 197301
rect 175779 197236 175780 197300
rect 175844 197236 175845 197300
rect 175779 197235 175845 197236
rect 175595 80204 175661 80205
rect 175595 80140 175596 80204
rect 175660 80140 175661 80204
rect 175595 80139 175661 80140
rect 175595 79932 175661 79933
rect 175595 79868 175596 79932
rect 175660 79868 175661 79932
rect 175595 79867 175661 79868
rect 175411 79524 175477 79525
rect 175411 79460 175412 79524
rect 175476 79460 175477 79524
rect 175411 79459 175477 79460
rect 175227 79252 175293 79253
rect 175227 79188 175228 79252
rect 175292 79188 175293 79252
rect 175227 79187 175293 79188
rect 175598 75581 175658 79867
rect 175782 79661 175842 197235
rect 175966 89730 176026 199003
rect 176334 195533 176394 199819
rect 182771 199748 182837 199749
rect 182771 199684 182772 199748
rect 182836 199684 182837 199748
rect 182771 199683 182837 199684
rect 180747 199612 180813 199613
rect 180747 199548 180748 199612
rect 180812 199548 180813 199612
rect 180747 199547 180813 199548
rect 176515 199476 176581 199477
rect 176515 199412 176516 199476
rect 176580 199412 176581 199476
rect 176515 199411 176581 199412
rect 176518 199069 176578 199411
rect 179643 199204 179709 199205
rect 179643 199140 179644 199204
rect 179708 199140 179709 199204
rect 179643 199139 179709 199140
rect 176515 199068 176581 199069
rect 176515 199004 176516 199068
rect 176580 199004 176581 199068
rect 176515 199003 176581 199004
rect 178355 198932 178421 198933
rect 178355 198868 178356 198932
rect 178420 198868 178421 198932
rect 178355 198867 178421 198868
rect 176699 198116 176765 198117
rect 176699 198052 176700 198116
rect 176764 198052 176765 198116
rect 176699 198051 176765 198052
rect 177067 198116 177133 198117
rect 177067 198052 177068 198116
rect 177132 198052 177133 198116
rect 177067 198051 177133 198052
rect 176702 197573 176762 198051
rect 176883 197980 176949 197981
rect 176883 197916 176884 197980
rect 176948 197916 176949 197980
rect 176883 197915 176949 197916
rect 176699 197572 176765 197573
rect 176699 197508 176700 197572
rect 176764 197508 176765 197572
rect 176699 197507 176765 197508
rect 176331 195532 176397 195533
rect 176331 195468 176332 195532
rect 176396 195468 176397 195532
rect 176331 195467 176397 195468
rect 175966 89670 176210 89730
rect 176150 79933 176210 89670
rect 176515 81292 176581 81293
rect 176515 81228 176516 81292
rect 176580 81228 176581 81292
rect 176515 81227 176581 81228
rect 176331 80612 176397 80613
rect 176331 80548 176332 80612
rect 176396 80548 176397 80612
rect 176331 80547 176397 80548
rect 176334 80205 176394 80547
rect 176331 80204 176397 80205
rect 176331 80140 176332 80204
rect 176396 80140 176397 80204
rect 176331 80139 176397 80140
rect 176147 79932 176213 79933
rect 176147 79868 176148 79932
rect 176212 79868 176213 79932
rect 176147 79867 176213 79868
rect 176331 79932 176397 79933
rect 176331 79868 176332 79932
rect 176396 79868 176397 79932
rect 176331 79867 176397 79868
rect 175963 79796 176029 79797
rect 175963 79732 175964 79796
rect 176028 79732 176029 79796
rect 175963 79731 176029 79732
rect 175779 79660 175845 79661
rect 175779 79596 175780 79660
rect 175844 79596 175845 79660
rect 175779 79595 175845 79596
rect 175966 79253 176026 79731
rect 175963 79252 176029 79253
rect 175963 79188 175964 79252
rect 176028 79188 176029 79252
rect 175963 79187 176029 79188
rect 176334 78434 176394 79867
rect 176518 78981 176578 81227
rect 176886 79797 176946 197915
rect 177070 79933 177130 198051
rect 177294 178954 177914 198000
rect 178171 197028 178237 197029
rect 178171 196964 178172 197028
rect 178236 196964 178237 197028
rect 178171 196963 178237 196964
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 177803 141268 177869 141269
rect 177803 141204 177804 141268
rect 177868 141204 177869 141268
rect 177803 141203 177869 141204
rect 177435 141132 177501 141133
rect 177435 141068 177436 141132
rect 177500 141068 177501 141132
rect 177435 141067 177501 141068
rect 177067 79932 177133 79933
rect 177067 79868 177068 79932
rect 177132 79868 177133 79932
rect 177438 79930 177498 141067
rect 177619 79932 177685 79933
rect 177619 79930 177620 79932
rect 177438 79870 177620 79930
rect 177067 79867 177133 79868
rect 177619 79868 177620 79870
rect 177684 79868 177685 79932
rect 177619 79867 177685 79868
rect 176883 79796 176949 79797
rect 176883 79732 176884 79796
rect 176948 79732 176949 79796
rect 176883 79731 176949 79732
rect 177070 79525 177130 79867
rect 177067 79524 177133 79525
rect 177067 79460 177068 79524
rect 177132 79460 177133 79524
rect 177067 79459 177133 79460
rect 176515 78980 176581 78981
rect 176515 78916 176516 78980
rect 176580 78916 176581 78980
rect 176515 78915 176581 78916
rect 177622 78573 177682 79867
rect 177806 79525 177866 141203
rect 177803 79524 177869 79525
rect 177803 79460 177804 79524
rect 177868 79460 177869 79524
rect 177803 79459 177869 79460
rect 177619 78572 177685 78573
rect 177619 78508 177620 78572
rect 177684 78508 177685 78572
rect 177619 78507 177685 78508
rect 176334 78374 176578 78434
rect 176331 78300 176397 78301
rect 176331 78236 176332 78300
rect 176396 78236 176397 78300
rect 176331 78235 176397 78236
rect 175963 78164 176029 78165
rect 175963 78100 175964 78164
rect 176028 78100 176029 78164
rect 175963 78099 176029 78100
rect 175595 75580 175661 75581
rect 175595 75516 175596 75580
rect 175660 75516 175661 75580
rect 175595 75515 175661 75516
rect 175966 70277 176026 78099
rect 176147 77212 176213 77213
rect 176147 77148 176148 77212
rect 176212 77148 176213 77212
rect 176147 77147 176213 77148
rect 175963 70276 176029 70277
rect 175963 70212 175964 70276
rect 176028 70212 176029 70276
rect 175963 70211 176029 70212
rect 176150 68781 176210 77147
rect 176147 68780 176213 68781
rect 176147 68716 176148 68780
rect 176212 68716 176213 68780
rect 176147 68715 176213 68716
rect 176334 60485 176394 78235
rect 176331 60484 176397 60485
rect 176331 60420 176332 60484
rect 176396 60420 176397 60484
rect 176331 60419 176397 60420
rect 175043 57220 175109 57221
rect 175043 57156 175044 57220
rect 175108 57156 175109 57220
rect 175043 57155 175109 57156
rect 176518 56133 176578 78374
rect 177067 77892 177133 77893
rect 177067 77828 177068 77892
rect 177132 77828 177133 77892
rect 177067 77827 177133 77828
rect 177070 74085 177130 77827
rect 177067 74084 177133 74085
rect 177067 74020 177068 74084
rect 177132 74020 177133 74084
rect 177067 74019 177133 74020
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 176515 56132 176581 56133
rect 176515 56068 176516 56132
rect 176580 56068 176581 56132
rect 176515 56067 176581 56068
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 70398
rect 178174 67285 178234 196963
rect 178358 70005 178418 198867
rect 179459 197708 179525 197709
rect 179459 197644 179460 197708
rect 179524 197644 179525 197708
rect 179459 197643 179525 197644
rect 178907 140044 178973 140045
rect 178907 139980 178908 140044
rect 178972 139980 178973 140044
rect 178907 139979 178973 139980
rect 178539 139772 178605 139773
rect 178539 139708 178540 139772
rect 178604 139708 178605 139772
rect 178539 139707 178605 139708
rect 178542 76805 178602 139707
rect 178910 77213 178970 139979
rect 179462 78981 179522 197643
rect 179646 80749 179706 199139
rect 180750 195990 180810 199547
rect 180931 197572 180997 197573
rect 180931 197508 180932 197572
rect 180996 197508 180997 197572
rect 180931 197507 180997 197508
rect 180566 195930 180810 195990
rect 180011 147116 180077 147117
rect 180011 147052 180012 147116
rect 180076 147052 180077 147116
rect 180011 147051 180077 147052
rect 179827 145756 179893 145757
rect 179827 145692 179828 145756
rect 179892 145692 179893 145756
rect 179827 145691 179893 145692
rect 179643 80748 179709 80749
rect 179643 80684 179644 80748
rect 179708 80684 179709 80748
rect 179643 80683 179709 80684
rect 179459 78980 179525 78981
rect 179459 78916 179460 78980
rect 179524 78916 179525 78980
rect 179459 78915 179525 78916
rect 178907 77212 178973 77213
rect 178907 77148 178908 77212
rect 178972 77148 178973 77212
rect 178907 77147 178973 77148
rect 178539 76804 178605 76805
rect 178539 76740 178540 76804
rect 178604 76740 178605 76804
rect 178539 76739 178605 76740
rect 179830 73677 179890 145691
rect 180014 77213 180074 147051
rect 180566 89730 180626 195930
rect 180566 89670 180810 89730
rect 180750 78981 180810 89670
rect 180934 79525 180994 197507
rect 181794 183454 182414 198000
rect 182587 195396 182653 195397
rect 182587 195332 182588 195396
rect 182652 195332 182653 195396
rect 182587 195331 182653 195332
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181115 150108 181181 150109
rect 181115 150044 181116 150108
rect 181180 150044 181181 150108
rect 181115 150043 181181 150044
rect 180931 79524 180997 79525
rect 180931 79460 180932 79524
rect 180996 79460 180997 79524
rect 180931 79459 180997 79460
rect 180747 78980 180813 78981
rect 180747 78916 180748 78980
rect 180812 78916 180813 78980
rect 180747 78915 180813 78916
rect 180011 77212 180077 77213
rect 180011 77148 180012 77212
rect 180076 77148 180077 77212
rect 180011 77147 180077 77148
rect 181118 75037 181178 150043
rect 181794 147454 182414 182898
rect 181299 147388 181365 147389
rect 181299 147324 181300 147388
rect 181364 147324 181365 147388
rect 181299 147323 181365 147324
rect 181115 75036 181181 75037
rect 181115 74972 181116 75036
rect 181180 74972 181181 75036
rect 181115 74971 181181 74972
rect 181302 73813 181362 147323
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181299 73812 181365 73813
rect 181299 73748 181300 73812
rect 181364 73748 181365 73812
rect 181299 73747 181365 73748
rect 179827 73676 179893 73677
rect 179827 73612 179828 73676
rect 179892 73612 179893 73676
rect 179827 73611 179893 73612
rect 178355 70004 178421 70005
rect 178355 69940 178356 70004
rect 178420 69940 178421 70004
rect 178355 69939 178421 69940
rect 178171 67284 178237 67285
rect 178171 67220 178172 67284
rect 178236 67220 178237 67284
rect 178171 67219 178237 67220
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 74898
rect 182590 53413 182650 195331
rect 182774 70141 182834 199683
rect 187003 198660 187069 198661
rect 187003 198596 187004 198660
rect 187068 198596 187069 198660
rect 187003 198595 187069 198596
rect 186294 187954 186914 198000
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186083 152692 186149 152693
rect 186083 152628 186084 152692
rect 186148 152628 186149 152692
rect 186083 152627 186149 152628
rect 185163 152556 185229 152557
rect 185163 152492 185164 152556
rect 185228 152492 185229 152556
rect 185163 152491 185229 152492
rect 182955 150244 183021 150245
rect 182955 150180 182956 150244
rect 183020 150180 183021 150244
rect 182955 150179 183021 150180
rect 182771 70140 182837 70141
rect 182771 70076 182772 70140
rect 182836 70076 182837 70140
rect 182771 70075 182837 70076
rect 182958 68917 183018 150179
rect 183139 149972 183205 149973
rect 183139 149908 183140 149972
rect 183204 149908 183205 149972
rect 183139 149907 183205 149908
rect 183142 72997 183202 149907
rect 183507 149836 183573 149837
rect 183507 149772 183508 149836
rect 183572 149772 183573 149836
rect 183507 149771 183573 149772
rect 183323 139500 183389 139501
rect 183323 139436 183324 139500
rect 183388 139436 183389 139500
rect 183323 139435 183389 139436
rect 183326 138957 183386 139435
rect 183323 138956 183389 138957
rect 183323 138892 183324 138956
rect 183388 138892 183389 138956
rect 183323 138891 183389 138892
rect 183510 74221 183570 149771
rect 184979 149700 185045 149701
rect 184979 149636 184980 149700
rect 185044 149636 185045 149700
rect 184979 149635 185045 149636
rect 183691 146980 183757 146981
rect 183691 146916 183692 146980
rect 183756 146916 183757 146980
rect 183691 146915 183757 146916
rect 183694 76397 183754 146915
rect 183875 141404 183941 141405
rect 183875 141340 183876 141404
rect 183940 141340 183941 141404
rect 183875 141339 183941 141340
rect 183878 93870 183938 141339
rect 184427 140452 184493 140453
rect 184427 140388 184428 140452
rect 184492 140388 184493 140452
rect 184427 140387 184493 140388
rect 184430 138413 184490 140387
rect 184427 138412 184493 138413
rect 184427 138348 184428 138412
rect 184492 138348 184493 138412
rect 184427 138347 184493 138348
rect 183878 93810 184122 93870
rect 183691 76396 183757 76397
rect 183691 76332 183692 76396
rect 183756 76332 183757 76396
rect 183691 76331 183757 76332
rect 183507 74220 183573 74221
rect 183507 74156 183508 74220
rect 183572 74156 183573 74220
rect 183507 74155 183573 74156
rect 183139 72996 183205 72997
rect 183139 72932 183140 72996
rect 183204 72932 183205 72996
rect 183139 72931 183205 72932
rect 184062 71501 184122 93810
rect 184982 71773 185042 149635
rect 185166 137869 185226 152491
rect 185347 152420 185413 152421
rect 185347 152356 185348 152420
rect 185412 152356 185413 152420
rect 185347 152355 185413 152356
rect 185350 138005 185410 152355
rect 185715 139772 185781 139773
rect 185715 139708 185716 139772
rect 185780 139708 185781 139772
rect 185715 139707 185781 139708
rect 185718 139093 185778 139707
rect 185715 139092 185781 139093
rect 185715 139028 185716 139092
rect 185780 139028 185781 139092
rect 185715 139027 185781 139028
rect 185347 138004 185413 138005
rect 185347 137940 185348 138004
rect 185412 137940 185413 138004
rect 185347 137939 185413 137940
rect 185163 137868 185229 137869
rect 185163 137804 185164 137868
rect 185228 137804 185229 137868
rect 185163 137803 185229 137804
rect 186086 127669 186146 152627
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 186267 138276 186333 138277
rect 186267 138212 186268 138276
rect 186332 138212 186333 138276
rect 186267 138211 186333 138212
rect 186083 127668 186149 127669
rect 186083 127604 186084 127668
rect 186148 127604 186149 127668
rect 186083 127603 186149 127604
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 186270 89730 186330 138211
rect 186086 89670 186330 89730
rect 186086 80070 186146 89670
rect 186086 80069 186330 80070
rect 186086 80068 186333 80069
rect 186086 80010 186268 80068
rect 186267 80004 186268 80010
rect 186332 80004 186333 80068
rect 186267 80003 186333 80004
rect 184979 71772 185045 71773
rect 184979 71708 184980 71772
rect 185044 71708 185045 71772
rect 184979 71707 185045 71708
rect 184059 71500 184125 71501
rect 184059 71436 184060 71500
rect 184124 71436 184125 71500
rect 184059 71435 184125 71436
rect 182955 68916 183021 68917
rect 182955 68852 182956 68916
rect 183020 68852 183021 68916
rect 182955 68851 183021 68852
rect 182587 53412 182653 53413
rect 182587 53348 182588 53412
rect 182652 53348 182653 53412
rect 182587 53347 182653 53348
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 187006 64701 187066 198595
rect 187190 143445 187250 212467
rect 187739 198524 187805 198525
rect 187739 198460 187740 198524
rect 187804 198460 187805 198524
rect 187739 198459 187805 198460
rect 187187 143444 187253 143445
rect 187187 143380 187188 143444
rect 187252 143380 187253 143444
rect 187187 143379 187253 143380
rect 187187 138140 187253 138141
rect 187187 138076 187188 138140
rect 187252 138076 187253 138140
rect 187187 138075 187253 138076
rect 187003 64700 187069 64701
rect 187003 64636 187004 64700
rect 187068 64636 187069 64700
rect 187003 64635 187069 64636
rect 187006 64293 187066 64635
rect 187003 64292 187069 64293
rect 187003 64228 187004 64292
rect 187068 64228 187069 64292
rect 187003 64227 187069 64228
rect 187190 62117 187250 138075
rect 187742 74085 187802 198459
rect 187923 197844 187989 197845
rect 187923 197780 187924 197844
rect 187988 197780 187989 197844
rect 187923 197779 187989 197780
rect 187926 78437 187986 197779
rect 189030 142901 189090 277475
rect 189211 276044 189277 276045
rect 189211 275980 189212 276044
rect 189276 275980 189277 276044
rect 189211 275979 189277 275980
rect 189027 142900 189093 142901
rect 189027 142836 189028 142900
rect 189092 142836 189093 142900
rect 189027 142835 189093 142836
rect 189214 142629 189274 275979
rect 190794 264454 191414 299898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 194547 265164 194613 265165
rect 194547 265100 194548 265164
rect 194612 265100 194613 265164
rect 194547 265099 194613 265100
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190499 262308 190565 262309
rect 190499 262244 190500 262308
rect 190564 262244 190565 262308
rect 190499 262243 190565 262244
rect 189579 260132 189645 260133
rect 189579 260068 189580 260132
rect 189644 260068 189645 260132
rect 189579 260067 189645 260068
rect 189395 198388 189461 198389
rect 189395 198324 189396 198388
rect 189460 198324 189461 198388
rect 189395 198323 189461 198324
rect 189211 142628 189277 142629
rect 189211 142564 189212 142628
rect 189276 142564 189277 142628
rect 189211 142563 189277 142564
rect 188291 140996 188357 140997
rect 188291 140932 188292 140996
rect 188356 140932 188357 140996
rect 188291 140931 188357 140932
rect 187923 78436 187989 78437
rect 187923 78372 187924 78436
rect 187988 78372 187989 78436
rect 187923 78371 187989 78372
rect 187926 77893 187986 78371
rect 187923 77892 187989 77893
rect 187923 77828 187924 77892
rect 187988 77828 187989 77892
rect 187923 77827 187989 77828
rect 187739 74084 187805 74085
rect 187739 74020 187740 74084
rect 187804 74020 187805 74084
rect 187739 74019 187805 74020
rect 187742 71229 187802 74019
rect 187739 71228 187805 71229
rect 187739 71164 187740 71228
rect 187804 71164 187805 71228
rect 187739 71163 187805 71164
rect 187187 62116 187253 62117
rect 187187 62052 187188 62116
rect 187252 62052 187253 62116
rect 187187 62051 187253 62052
rect 188294 59397 188354 140931
rect 188475 140180 188541 140181
rect 188475 140116 188476 140180
rect 188540 140116 188541 140180
rect 188475 140115 188541 140116
rect 188478 125629 188538 140115
rect 189027 139772 189093 139773
rect 189027 139708 189028 139772
rect 189092 139708 189093 139772
rect 189027 139707 189093 139708
rect 188475 125628 188541 125629
rect 188475 125564 188476 125628
rect 188540 125564 188541 125628
rect 188475 125563 188541 125564
rect 189030 75037 189090 139707
rect 189027 75036 189093 75037
rect 189027 74972 189028 75036
rect 189092 74972 189093 75036
rect 189027 74971 189093 74972
rect 189030 67557 189090 74971
rect 189027 67556 189093 67557
rect 189027 67492 189028 67556
rect 189092 67492 189093 67556
rect 189027 67491 189093 67492
rect 189398 65789 189458 198323
rect 189582 142765 189642 260067
rect 190502 144261 190562 262243
rect 190794 262000 191414 263898
rect 193443 262716 193509 262717
rect 193443 262652 193444 262716
rect 193508 262652 193509 262716
rect 193443 262651 193509 262652
rect 191971 262580 192037 262581
rect 191971 262516 191972 262580
rect 192036 262516 192037 262580
rect 191971 262515 192037 262516
rect 191787 259724 191853 259725
rect 191787 259660 191788 259724
rect 191852 259660 191853 259724
rect 191787 259659 191853 259660
rect 190794 192454 191414 198000
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190499 144260 190565 144261
rect 190499 144196 190500 144260
rect 190564 144196 190565 144260
rect 190499 144195 190565 144196
rect 189579 142764 189645 142765
rect 189579 142700 189580 142764
rect 189644 142700 189645 142764
rect 189579 142699 189645 142700
rect 190794 142000 191414 155898
rect 191790 142085 191850 259659
rect 191974 143989 192034 262515
rect 192155 262308 192221 262309
rect 192155 262244 192156 262308
rect 192220 262244 192221 262308
rect 192155 262243 192221 262244
rect 192158 144125 192218 262243
rect 193259 197164 193325 197165
rect 193259 197100 193260 197164
rect 193324 197100 193325 197164
rect 193259 197099 193325 197100
rect 192523 146164 192589 146165
rect 192523 146100 192524 146164
rect 192588 146100 192589 146164
rect 192523 146099 192589 146100
rect 192155 144124 192221 144125
rect 192155 144060 192156 144124
rect 192220 144060 192221 144124
rect 192155 144059 192221 144060
rect 191971 143988 192037 143989
rect 191971 143924 191972 143988
rect 192036 143924 192037 143988
rect 191971 143923 192037 143924
rect 191787 142084 191853 142085
rect 191787 142020 191788 142084
rect 191852 142020 191853 142084
rect 191787 142019 191853 142020
rect 190499 141540 190565 141541
rect 190499 141476 190500 141540
rect 190564 141476 190565 141540
rect 190499 141475 190565 141476
rect 189579 139908 189645 139909
rect 189579 139844 189580 139908
rect 189644 139844 189645 139908
rect 189579 139843 189645 139844
rect 189582 111893 189642 139843
rect 189579 111892 189645 111893
rect 189579 111828 189580 111892
rect 189644 111828 189645 111892
rect 189579 111827 189645 111828
rect 189395 65788 189461 65789
rect 189395 65724 189396 65788
rect 189460 65724 189461 65788
rect 189395 65723 189461 65724
rect 188291 59396 188357 59397
rect 188291 59332 188292 59396
rect 188356 59332 188357 59396
rect 188291 59331 188357 59332
rect 190502 49061 190562 141475
rect 192339 140860 192405 140861
rect 192339 140796 192340 140860
rect 192404 140796 192405 140860
rect 192339 140795 192405 140796
rect 190867 140724 190933 140725
rect 190867 140660 190868 140724
rect 190932 140660 190933 140724
rect 190867 140659 190933 140660
rect 190870 79253 190930 140659
rect 191603 140316 191669 140317
rect 191603 140252 191604 140316
rect 191668 140252 191669 140316
rect 191603 140251 191669 140252
rect 190867 79252 190933 79253
rect 190867 79188 190868 79252
rect 190932 79188 190933 79252
rect 190867 79187 190933 79188
rect 190499 49060 190565 49061
rect 190499 48996 190500 49060
rect 190564 48996 190565 49060
rect 190499 48995 190565 48996
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 78000
rect 191606 76669 191666 140251
rect 191971 139908 192037 139909
rect 191971 139844 191972 139908
rect 192036 139844 192037 139908
rect 191971 139843 192037 139844
rect 191974 77077 192034 139843
rect 191971 77076 192037 77077
rect 191971 77012 191972 77076
rect 192036 77012 192037 77076
rect 191971 77011 192037 77012
rect 191603 76668 191669 76669
rect 191603 76604 191604 76668
rect 191668 76604 191669 76668
rect 191603 76603 191669 76604
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 192342 45661 192402 140795
rect 192526 73949 192586 146099
rect 193262 75581 193322 197099
rect 193446 144397 193506 262651
rect 193627 262444 193693 262445
rect 193627 262380 193628 262444
rect 193692 262380 193693 262444
rect 193627 262379 193693 262380
rect 193630 144941 193690 262379
rect 193811 147660 193877 147661
rect 193811 147596 193812 147660
rect 193876 147596 193877 147660
rect 193811 147595 193877 147596
rect 193627 144940 193693 144941
rect 193627 144876 193628 144940
rect 193692 144876 193693 144940
rect 193627 144875 193693 144876
rect 193443 144396 193509 144397
rect 193443 144332 193444 144396
rect 193508 144332 193509 144396
rect 193443 144331 193509 144332
rect 193259 75580 193325 75581
rect 193259 75516 193260 75580
rect 193324 75516 193325 75580
rect 193259 75515 193325 75516
rect 193814 74357 193874 147595
rect 193995 146028 194061 146029
rect 193995 145964 193996 146028
rect 194060 145964 194061 146028
rect 193995 145963 194061 145964
rect 193998 79389 194058 145963
rect 194550 144533 194610 265099
rect 195294 232954 195914 268398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 197491 265436 197557 265437
rect 197491 265372 197492 265436
rect 197556 265372 197557 265436
rect 197491 265371 197557 265372
rect 196203 265300 196269 265301
rect 196203 265236 196204 265300
rect 196268 265236 196269 265300
rect 196203 265235 196269 265236
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 196019 195124 196085 195125
rect 196019 195060 196020 195124
rect 196084 195060 196085 195124
rect 196019 195059 196085 195060
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195099 146980 195165 146981
rect 195099 146916 195100 146980
rect 195164 146916 195165 146980
rect 195099 146915 195165 146916
rect 194547 144532 194613 144533
rect 194547 144468 194548 144532
rect 194612 144468 194613 144532
rect 194547 144467 194613 144468
rect 193995 79388 194061 79389
rect 193995 79324 193996 79388
rect 194060 79324 194061 79388
rect 193995 79323 194061 79324
rect 193811 74356 193877 74357
rect 193811 74292 193812 74356
rect 193876 74292 193877 74356
rect 193811 74291 193877 74292
rect 192523 73948 192589 73949
rect 192523 73884 192524 73948
rect 192588 73884 192589 73948
rect 192523 73883 192589 73884
rect 195102 65517 195162 146915
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 195099 65516 195165 65517
rect 195099 65452 195100 65516
rect 195164 65452 195165 65516
rect 195099 65451 195165 65452
rect 195294 52954 195914 88398
rect 196022 62117 196082 195059
rect 196206 144669 196266 265235
rect 197307 195804 197373 195805
rect 197307 195740 197308 195804
rect 197372 195740 197373 195804
rect 197307 195739 197373 195740
rect 196387 147524 196453 147525
rect 196387 147460 196388 147524
rect 196452 147460 196453 147524
rect 196387 147459 196453 147460
rect 196203 144668 196269 144669
rect 196203 144604 196204 144668
rect 196268 144604 196269 144668
rect 196203 144603 196269 144604
rect 196390 75445 196450 147459
rect 196571 145892 196637 145893
rect 196571 145828 196572 145892
rect 196636 145828 196637 145892
rect 196571 145827 196637 145828
rect 196387 75444 196453 75445
rect 196387 75380 196388 75444
rect 196452 75380 196453 75444
rect 196387 75379 196453 75380
rect 196574 72861 196634 145827
rect 196571 72860 196637 72861
rect 196571 72796 196572 72860
rect 196636 72796 196637 72860
rect 196571 72795 196637 72796
rect 197310 62933 197370 195739
rect 197494 144805 197554 265371
rect 197675 265028 197741 265029
rect 197675 264964 197676 265028
rect 197740 264964 197741 265028
rect 197675 264963 197741 264964
rect 197678 145621 197738 264963
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199331 198796 199397 198797
rect 199331 198732 199332 198796
rect 199396 198732 199397 198796
rect 199331 198731 199397 198732
rect 198963 198252 199029 198253
rect 198963 198188 198964 198252
rect 199028 198188 199029 198252
rect 198963 198187 199029 198188
rect 198779 195940 198845 195941
rect 198779 195876 198780 195940
rect 198844 195876 198845 195940
rect 198779 195875 198845 195876
rect 198043 147252 198109 147253
rect 198043 147188 198044 147252
rect 198108 147188 198109 147252
rect 198043 147187 198109 147188
rect 197859 146300 197925 146301
rect 197859 146236 197860 146300
rect 197924 146236 197925 146300
rect 197859 146235 197925 146236
rect 197675 145620 197741 145621
rect 197675 145556 197676 145620
rect 197740 145556 197741 145620
rect 197675 145555 197741 145556
rect 197491 144804 197557 144805
rect 197491 144740 197492 144804
rect 197556 144740 197557 144804
rect 197491 144739 197557 144740
rect 197491 71636 197557 71637
rect 197491 71572 197492 71636
rect 197556 71572 197557 71636
rect 197491 71571 197557 71572
rect 197494 71093 197554 71571
rect 197491 71092 197557 71093
rect 197491 71028 197492 71092
rect 197556 71028 197557 71092
rect 197491 71027 197557 71028
rect 197862 64837 197922 146235
rect 198046 71093 198106 147187
rect 198043 71092 198109 71093
rect 198043 71028 198044 71092
rect 198108 71028 198109 71092
rect 198043 71027 198109 71028
rect 198782 68917 198842 195875
rect 198966 80749 199026 198187
rect 198963 80748 199029 80749
rect 198963 80684 198964 80748
rect 199028 80684 199029 80748
rect 198963 80683 199029 80684
rect 199334 78981 199394 198731
rect 199794 165454 200414 200898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 200619 195668 200685 195669
rect 200619 195604 200620 195668
rect 200684 195604 200685 195668
rect 200619 195603 200685 195604
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 198963 78980 199029 78981
rect 198963 78916 198964 78980
rect 199028 78916 199029 78980
rect 198963 78915 199029 78916
rect 199331 78980 199397 78981
rect 199331 78916 199332 78980
rect 199396 78916 199397 78980
rect 199331 78915 199397 78916
rect 198966 78165 199026 78915
rect 198963 78164 199029 78165
rect 198963 78100 198964 78164
rect 199028 78100 199029 78164
rect 198963 78099 199029 78100
rect 198779 68916 198845 68917
rect 198779 68852 198780 68916
rect 198844 68852 198845 68916
rect 198779 68851 198845 68852
rect 197859 64836 197925 64837
rect 197859 64772 197860 64836
rect 197924 64772 197925 64836
rect 197859 64771 197925 64772
rect 197862 64157 197922 64771
rect 197859 64156 197925 64157
rect 197859 64092 197860 64156
rect 197924 64092 197925 64156
rect 197859 64091 197925 64092
rect 197307 62932 197373 62933
rect 197307 62868 197308 62932
rect 197372 62868 197373 62932
rect 197307 62867 197373 62868
rect 196019 62116 196085 62117
rect 196019 62052 196020 62116
rect 196084 62052 196085 62116
rect 196019 62051 196085 62052
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 192339 45660 192405 45661
rect 192339 45596 192340 45660
rect 192404 45596 192405 45660
rect 192339 45595 192405 45596
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 200622 56133 200682 195603
rect 200987 195532 201053 195533
rect 200987 195468 200988 195532
rect 201052 195468 201053 195532
rect 200987 195467 201053 195468
rect 200803 195260 200869 195261
rect 200803 195196 200804 195260
rect 200868 195196 200869 195260
rect 200803 195195 200869 195196
rect 200806 57221 200866 195195
rect 200990 59941 201050 195467
rect 201723 194036 201789 194037
rect 201723 193972 201724 194036
rect 201788 193972 201789 194036
rect 201723 193971 201789 193972
rect 201539 193900 201605 193901
rect 201539 193836 201540 193900
rect 201604 193836 201605 193900
rect 201539 193835 201605 193836
rect 201171 147796 201237 147797
rect 201171 147732 201172 147796
rect 201236 147732 201237 147796
rect 201171 147731 201237 147732
rect 201174 74550 201234 147731
rect 201174 74490 201418 74550
rect 201358 70277 201418 74490
rect 201355 70276 201421 70277
rect 201355 70212 201356 70276
rect 201420 70212 201421 70276
rect 201355 70211 201421 70212
rect 201358 69597 201418 70211
rect 201355 69596 201421 69597
rect 201355 69532 201356 69596
rect 201420 69532 201421 69596
rect 201355 69531 201421 69532
rect 200987 59940 201053 59941
rect 200987 59876 200988 59940
rect 201052 59876 201053 59940
rect 200987 59875 201053 59876
rect 200803 57220 200869 57221
rect 200803 57156 200804 57220
rect 200868 57156 200869 57220
rect 200803 57155 200869 57156
rect 200619 56132 200685 56133
rect 200619 56068 200620 56132
rect 200684 56068 200685 56132
rect 200619 56067 200685 56068
rect 201355 56132 201421 56133
rect 201355 56068 201356 56132
rect 201420 56068 201421 56132
rect 201355 56067 201421 56068
rect 201358 55861 201418 56067
rect 201355 55860 201421 55861
rect 201355 55796 201356 55860
rect 201420 55796 201421 55860
rect 201355 55795 201421 55796
rect 201542 46205 201602 193835
rect 201726 55181 201786 193971
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 203011 150380 203077 150381
rect 203011 150316 203012 150380
rect 203076 150316 203077 150380
rect 203011 150315 203077 150316
rect 201723 55180 201789 55181
rect 201723 55116 201724 55180
rect 201788 55116 201789 55180
rect 201723 55115 201789 55116
rect 203014 50965 203074 150315
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 203011 50964 203077 50965
rect 203011 50900 203012 50964
rect 203076 50900 203077 50964
rect 203011 50899 203077 50900
rect 201539 46204 201605 46205
rect 201539 46140 201540 46204
rect 201604 46140 201605 46204
rect 201539 46139 201605 46140
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 124250 255218 124486 255454
rect 124250 254898 124486 255134
rect 154970 255218 155206 255454
rect 154970 254898 155206 255134
rect 185690 255218 185926 255454
rect 185690 254898 185926 255134
rect 139610 223718 139846 223954
rect 139610 223398 139846 223634
rect 170330 223718 170566 223954
rect 170330 223398 170566 223634
rect 124250 219218 124486 219454
rect 124250 218898 124486 219134
rect 154970 219218 155206 219454
rect 154970 218898 155206 219134
rect 185690 219218 185926 219454
rect 185690 218898 185926 219134
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 124250 255454
rect 124486 255218 154970 255454
rect 155206 255218 185690 255454
rect 185926 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 124250 255134
rect 124486 254898 154970 255134
rect 155206 254898 185690 255134
rect 185926 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 139610 223954
rect 139846 223718 170330 223954
rect 170566 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 139610 223634
rect 139846 223398 170330 223634
rect 170566 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 124250 219454
rect 124486 219218 154970 219454
rect 155206 219218 185690 219454
rect 185926 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 124250 219134
rect 124486 218898 154970 219134
rect 155206 218898 185690 219134
rect 185926 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use pixel_macro  pixel_macro0
timestamp 0
transform 1 0 120000 0 1 200000
box 1066 0 68854 60000
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 1066 0 68854 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 262000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 198000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 262000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 262000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 262000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 142000 191414 198000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 262000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 262000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 262000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 262000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 262000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 262000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 262000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 262000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 198000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 262000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 262000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 198000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 262000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 262000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 198000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 262000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
