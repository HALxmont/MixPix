magic
tech sky130B
magscale 1 2
timestamp 1668044308
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 207658 700680 207664 700732
rect 207716 700720 207722 700732
rect 218974 700720 218980 700732
rect 207716 700692 218980 700720
rect 207716 700680 207722 700692
rect 218974 700680 218980 700692
rect 219032 700680 219038 700732
rect 192478 700612 192484 700664
rect 192536 700652 192542 700664
rect 267642 700652 267648 700664
rect 192536 700624 267648 700652
rect 192536 700612 192542 700624
rect 267642 700612 267648 700624
rect 267700 700612 267706 700664
rect 206278 700544 206284 700596
rect 206336 700584 206342 700596
rect 283834 700584 283840 700596
rect 206336 700556 283840 700584
rect 206336 700544 206342 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 203518 700476 203524 700528
rect 203576 700516 203582 700528
rect 348786 700516 348792 700528
rect 203576 700488 348792 700516
rect 203576 700476 203582 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 200758 700408 200764 700460
rect 200816 700448 200822 700460
rect 413646 700448 413652 700460
rect 200816 700420 413652 700448
rect 200816 700408 200822 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 199378 700340 199384 700392
rect 199436 700380 199442 700392
rect 478506 700380 478512 700392
rect 199436 700352 478512 700380
rect 199436 700340 199442 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 137830 700272 137836 700324
rect 137888 700312 137894 700324
rect 190454 700312 190460 700324
rect 137888 700284 190460 700312
rect 137888 700272 137894 700284
rect 190454 700272 190460 700284
rect 190512 700272 190518 700324
rect 197998 700272 198004 700324
rect 198056 700312 198062 700324
rect 543458 700312 543464 700324
rect 198056 700284 543464 700312
rect 198056 700272 198062 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106918 699700 106924 699712
rect 105504 699672 106924 699700
rect 105504 699660 105510 699672
rect 106918 699660 106924 699672
rect 106976 699660 106982 699712
rect 193858 699660 193864 699712
rect 193916 699700 193922 699712
rect 202782 699700 202788 699712
rect 193916 699672 202788 699700
rect 193916 699660 193922 699672
rect 202782 699660 202788 699672
rect 202840 699660 202846 699712
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 196618 683136 196624 683188
rect 196676 683176 196682 683188
rect 580166 683176 580172 683188
rect 196676 683148 580172 683176
rect 196676 683136 196682 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 116578 656928 116584 656940
rect 3476 656900 116584 656928
rect 3476 656888 3482 656900
rect 116578 656888 116584 656900
rect 116636 656888 116642 656940
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 7558 632108 7564 632120
rect 3476 632080 7564 632108
rect 3476 632068 3482 632080
rect 7558 632068 7564 632080
rect 7616 632068 7622 632120
rect 193950 630640 193956 630692
rect 194008 630680 194014 630692
rect 580166 630680 580172 630692
rect 194008 630652 580172 630680
rect 194008 630640 194014 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 120718 616836 120724 616888
rect 120776 616876 120782 616888
rect 580166 616876 580172 616888
rect 120776 616848 580172 616876
rect 120776 616836 120782 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 17218 579680 17224 579692
rect 3384 579652 17224 579680
rect 3384 579640 3390 579652
rect 17218 579640 17224 579652
rect 17276 579640 17282 579692
rect 194042 576852 194048 576904
rect 194100 576892 194106 576904
rect 579614 576892 579620 576904
rect 194100 576864 579620 576892
rect 194100 576852 194106 576864
rect 579614 576852 579620 576864
rect 579672 576852 579678 576904
rect 120810 563048 120816 563100
rect 120868 563088 120874 563100
rect 580166 563088 580172 563100
rect 120868 563060 580172 563088
rect 120868 563048 120874 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 116670 553432 116676 553444
rect 3384 553404 116676 553432
rect 3384 553392 3390 553404
rect 116670 553392 116676 553404
rect 116728 553392 116734 553444
rect 3326 527824 3332 527876
rect 3384 527864 3390 527876
rect 8938 527864 8944 527876
rect 3384 527836 8944 527864
rect 3384 527824 3390 527836
rect 8938 527824 8944 527836
rect 8996 527824 9002 527876
rect 194134 524424 194140 524476
rect 194192 524464 194198 524476
rect 579798 524464 579804 524476
rect 194192 524436 579804 524464
rect 194192 524424 194198 524436
rect 579798 524424 579804 524436
rect 579856 524424 579862 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 190546 514808 190552 514820
rect 3384 514780 190552 514808
rect 3384 514768 3390 514780
rect 190546 514768 190552 514780
rect 190604 514768 190610 514820
rect 120902 510620 120908 510672
rect 120960 510660 120966 510672
rect 579982 510660 579988 510672
rect 120960 510632 579988 510660
rect 120960 510620 120966 510632
rect 579982 510620 579988 510632
rect 580040 510620 580046 510672
rect 118694 485052 118700 485104
rect 118752 485092 118758 485104
rect 580534 485092 580540 485104
rect 118752 485064 580540 485092
rect 118752 485052 118758 485064
rect 580534 485052 580540 485064
rect 580592 485052 580598 485104
rect 221458 470568 221464 470620
rect 221516 470608 221522 470620
rect 579614 470608 579620 470620
rect 221516 470580 579620 470608
rect 221516 470568 221522 470580
rect 579614 470568 579620 470580
rect 579672 470568 579678 470620
rect 3050 462340 3056 462392
rect 3108 462380 3114 462392
rect 189718 462380 189724 462392
rect 3108 462352 189724 462380
rect 3108 462340 3114 462352
rect 189718 462340 189724 462352
rect 189776 462340 189782 462392
rect 3878 461592 3884 461644
rect 3936 461632 3942 461644
rect 48958 461632 48964 461644
rect 3936 461604 48964 461632
rect 3936 461592 3942 461604
rect 48958 461592 48964 461604
rect 49016 461592 49022 461644
rect 120994 456764 121000 456816
rect 121052 456804 121058 456816
rect 579614 456804 579620 456816
rect 121052 456776 579620 456804
rect 121052 456764 121058 456776
rect 579614 456764 579620 456776
rect 579672 456764 579678 456816
rect 2958 448536 2964 448588
rect 3016 448576 3022 448588
rect 84838 448576 84844 448588
rect 3016 448548 84844 448576
rect 3016 448536 3022 448548
rect 84838 448536 84844 448548
rect 84896 448536 84902 448588
rect 3326 422288 3332 422340
rect 3384 422328 3390 422340
rect 10318 422328 10324 422340
rect 3384 422300 10324 422328
rect 3384 422288 3390 422300
rect 10318 422288 10324 422300
rect 10376 422288 10382 422340
rect 192570 418140 192576 418192
rect 192628 418180 192634 418192
rect 579706 418180 579712 418192
rect 192628 418152 579712 418180
rect 192628 418140 192634 418152
rect 579706 418140 579712 418152
rect 579764 418140 579770 418192
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 189074 409884 189080 409896
rect 3384 409856 189080 409884
rect 3384 409844 3390 409856
rect 189074 409844 189080 409856
rect 189132 409844 189138 409896
rect 118602 404336 118608 404388
rect 118660 404376 118666 404388
rect 580166 404376 580172 404388
rect 118660 404348 580172 404376
rect 118660 404336 118666 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 112438 397508 112444 397520
rect 3384 397480 112444 397508
rect 3384 397468 3390 397480
rect 112438 397468 112444 397480
rect 112496 397468 112502 397520
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 84930 371260 84936 371272
rect 3384 371232 84936 371260
rect 3384 371220 3390 371232
rect 84930 371220 84936 371232
rect 84988 371220 84994 371272
rect 360838 364352 360844 364404
rect 360896 364392 360902 364404
rect 580166 364392 580172 364404
rect 360896 364364 580172 364392
rect 360896 364352 360902 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 118510 351908 118516 351960
rect 118568 351948 118574 351960
rect 580166 351948 580172 351960
rect 118568 351920 580172 351948
rect 118568 351908 118574 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 121086 345080 121092 345092
rect 3384 345052 121092 345080
rect 3384 345040 3390 345052
rect 121086 345040 121092 345052
rect 121144 345040 121150 345092
rect 3142 318792 3148 318844
rect 3200 318832 3206 318844
rect 13078 318832 13084 318844
rect 3200 318804 13084 318832
rect 3200 318792 3206 318804
rect 13078 318792 13084 318804
rect 13136 318792 13142 318844
rect 359458 311856 359464 311908
rect 359516 311896 359522 311908
rect 580166 311896 580172 311908
rect 359516 311868 580172 311896
rect 359516 311856 359522 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 3326 304988 3332 305040
rect 3384 305028 3390 305040
rect 185578 305028 185584 305040
rect 3384 305000 185584 305028
rect 3384 304988 3390 305000
rect 185578 304988 185584 305000
rect 185636 304988 185642 305040
rect 146938 298120 146944 298172
rect 146996 298160 147002 298172
rect 580166 298160 580172 298172
rect 146996 298132 580172 298160
rect 146996 298120 147002 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3234 266364 3240 266416
rect 3292 266404 3298 266416
rect 18598 266404 18604 266416
rect 3292 266376 18604 266404
rect 3292 266364 3298 266376
rect 18598 266364 18604 266376
rect 18656 266364 18662 266416
rect 202138 258068 202144 258120
rect 202196 258108 202202 258120
rect 580166 258108 580172 258120
rect 202196 258080 580172 258108
rect 202196 258068 202202 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 2866 253920 2872 253972
rect 2924 253960 2930 253972
rect 190638 253960 190644 253972
rect 2924 253932 190644 253960
rect 2924 253920 2930 253932
rect 190638 253920 190644 253932
rect 190696 253920 190702 253972
rect 122098 244264 122104 244316
rect 122156 244304 122162 244316
rect 580166 244304 580172 244316
rect 122156 244276 580172 244304
rect 122156 244264 122162 244276
rect 580166 244264 580172 244276
rect 580224 244264 580230 244316
rect 194226 231820 194232 231872
rect 194284 231860 194290 231872
rect 579798 231860 579804 231872
rect 194284 231832 579804 231860
rect 194284 231820 194290 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 225598 218016 225604 218068
rect 225656 218056 225662 218068
rect 579982 218056 579988 218068
rect 225656 218028 579988 218056
rect 225656 218016 225662 218028
rect 579982 218016 579988 218028
rect 580040 218016 580046 218068
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 31018 213976 31024 213988
rect 3384 213948 31024 213976
rect 3384 213936 3390 213948
rect 31018 213936 31024 213948
rect 31076 213936 31082 213988
rect 147030 205640 147036 205692
rect 147088 205680 147094 205692
rect 580166 205680 580172 205692
rect 147088 205652 580172 205680
rect 147088 205640 147094 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 3326 201492 3332 201544
rect 3384 201532 3390 201544
rect 189258 201532 189264 201544
rect 3384 201504 189264 201532
rect 3384 201492 3390 201504
rect 189258 201492 189264 201504
rect 189316 201492 189322 201544
rect 192662 191836 192668 191888
rect 192720 191876 192726 191888
rect 580166 191876 580172 191888
rect 192720 191848 580172 191876
rect 192720 191836 192726 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 3326 187688 3332 187740
rect 3384 187728 3390 187740
rect 119338 187728 119344 187740
rect 3384 187700 119344 187728
rect 3384 187688 3390 187700
rect 119338 187688 119344 187700
rect 119396 187688 119402 187740
rect 224218 178032 224224 178084
rect 224276 178072 224282 178084
rect 580166 178072 580172 178084
rect 224276 178044 580172 178072
rect 224276 178032 224282 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 122190 165588 122196 165640
rect 122248 165628 122254 165640
rect 580166 165628 580172 165640
rect 122248 165600 580172 165628
rect 122248 165588 122254 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 3326 162868 3332 162920
rect 3384 162908 3390 162920
rect 14458 162908 14464 162920
rect 3384 162880 14464 162908
rect 3384 162868 3390 162880
rect 14458 162868 14464 162880
rect 14516 162868 14522 162920
rect 3786 160692 3792 160744
rect 3844 160732 3850 160744
rect 189350 160732 189356 160744
rect 3844 160704 189356 160732
rect 3844 160692 3850 160704
rect 189350 160692 189356 160704
rect 189408 160692 189414 160744
rect 192754 151784 192760 151836
rect 192812 151824 192818 151836
rect 579982 151824 579988 151836
rect 192812 151796 579988 151824
rect 192812 151784 192818 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 3510 149880 3516 149932
rect 3568 149920 3574 149932
rect 3786 149920 3792 149932
rect 3568 149892 3792 149920
rect 3568 149880 3574 149892
rect 3786 149880 3792 149892
rect 3844 149880 3850 149932
rect 3510 148316 3516 148368
rect 3568 148356 3574 148368
rect 191190 148356 191196 148368
rect 3568 148328 191196 148356
rect 3568 148316 3574 148328
rect 191190 148316 191196 148328
rect 191248 148316 191254 148368
rect 119246 146956 119252 147008
rect 119304 146996 119310 147008
rect 234614 146996 234620 147008
rect 119304 146968 234620 146996
rect 119304 146956 119310 146968
rect 234614 146956 234620 146968
rect 234672 146956 234678 147008
rect 3602 146888 3608 146940
rect 3660 146928 3666 146940
rect 190822 146928 190828 146940
rect 3660 146900 190828 146928
rect 3660 146888 3666 146900
rect 190822 146888 190828 146900
rect 190880 146888 190886 146940
rect 118970 145596 118976 145648
rect 119028 145636 119034 145648
rect 299474 145636 299480 145648
rect 119028 145608 299480 145636
rect 119028 145596 119034 145608
rect 299474 145596 299480 145608
rect 299532 145596 299538 145648
rect 3786 145528 3792 145580
rect 3844 145568 3850 145580
rect 189442 145568 189448 145580
rect 3844 145540 189448 145568
rect 3844 145528 3850 145540
rect 189442 145528 189448 145540
rect 189500 145528 189506 145580
rect 23474 144236 23480 144288
rect 23532 144276 23538 144288
rect 189534 144276 189540 144288
rect 23532 144248 189540 144276
rect 23532 144236 23538 144248
rect 189534 144236 189540 144248
rect 189592 144236 189598 144288
rect 119062 144168 119068 144220
rect 119120 144208 119126 144220
rect 364334 144208 364340 144220
rect 119120 144180 364340 144208
rect 119120 144168 119126 144180
rect 364334 144168 364340 144180
rect 364392 144168 364398 144220
rect 118234 142944 118240 142996
rect 118292 142984 118298 142996
rect 146938 142984 146944 142996
rect 118292 142956 146944 142984
rect 118292 142944 118298 142956
rect 146938 142944 146944 142956
rect 146996 142944 147002 142996
rect 3878 142876 3884 142928
rect 3936 142916 3942 142928
rect 191098 142916 191104 142928
rect 3936 142888 191104 142916
rect 3936 142876 3942 142888
rect 191098 142876 191104 142888
rect 191156 142876 191162 142928
rect 119154 142808 119160 142860
rect 119212 142848 119218 142860
rect 429194 142848 429200 142860
rect 119212 142820 429200 142848
rect 119212 142808 119218 142820
rect 429194 142808 429200 142820
rect 429252 142808 429258 142860
rect 118418 141516 118424 141568
rect 118476 141556 118482 141568
rect 147030 141556 147036 141568
rect 118476 141528 147036 141556
rect 118476 141516 118482 141528
rect 147030 141516 147036 141528
rect 147088 141516 147094 141568
rect 88334 141448 88340 141500
rect 88392 141488 88398 141500
rect 191006 141488 191012 141500
rect 88392 141460 191012 141488
rect 88392 141448 88398 141460
rect 191006 141448 191012 141460
rect 191064 141448 191070 141500
rect 118878 141380 118884 141432
rect 118936 141420 118942 141432
rect 494054 141420 494060 141432
rect 118936 141392 494060 141420
rect 118936 141380 118942 141392
rect 494054 141380 494060 141392
rect 494112 141380 494118 141432
rect 185578 140496 185584 140548
rect 185636 140536 185642 140548
rect 192018 140536 192024 140548
rect 185636 140508 192024 140536
rect 185636 140496 185642 140508
rect 192018 140496 192024 140508
rect 192076 140496 192082 140548
rect 153194 140156 153200 140208
rect 153252 140196 153258 140208
rect 190914 140196 190920 140208
rect 153252 140168 190920 140196
rect 153252 140156 153258 140168
rect 190914 140156 190920 140168
rect 190972 140156 190978 140208
rect 118050 140088 118056 140140
rect 118108 140128 118114 140140
rect 169754 140128 169760 140140
rect 118108 140100 169760 140128
rect 118108 140088 118114 140100
rect 169754 140088 169760 140100
rect 169812 140088 169818 140140
rect 118786 140020 118792 140072
rect 118844 140060 118850 140072
rect 558914 140060 558920 140072
rect 118844 140032 558920 140060
rect 118844 140020 118850 140032
rect 558914 140020 558920 140032
rect 558972 140020 558978 140072
rect 118142 139544 118148 139596
rect 118200 139584 118206 139596
rect 122098 139584 122104 139596
rect 118200 139556 122104 139584
rect 118200 139544 118206 139556
rect 122098 139544 122104 139556
rect 122156 139544 122162 139596
rect 118326 139476 118332 139528
rect 118384 139516 118390 139528
rect 122190 139516 122196 139528
rect 118384 139488 122196 139516
rect 118384 139476 118390 139488
rect 122190 139476 122196 139488
rect 122248 139476 122254 139528
rect 3602 139408 3608 139460
rect 3660 139448 3666 139460
rect 191926 139448 191932 139460
rect 3660 139420 191932 139448
rect 3660 139408 3666 139420
rect 191926 139408 191932 139420
rect 191984 139408 191990 139460
rect 7650 136688 7656 136740
rect 7708 136728 7714 136740
rect 117314 136728 117320 136740
rect 7708 136700 117320 136728
rect 7708 136688 7714 136700
rect 117314 136688 117320 136700
rect 117372 136688 117378 136740
rect 3510 136620 3516 136672
rect 3568 136660 3574 136672
rect 119430 136660 119436 136672
rect 3568 136632 119436 136660
rect 3568 136620 3574 136632
rect 119430 136620 119436 136632
rect 119488 136620 119494 136672
rect 9030 135260 9036 135312
rect 9088 135300 9094 135312
rect 117314 135300 117320 135312
rect 9088 135272 117320 135300
rect 9088 135260 9094 135272
rect 117314 135260 117320 135272
rect 117372 135260 117378 135312
rect 21358 133900 21364 133952
rect 21416 133940 21422 133952
rect 117314 133940 117320 133952
rect 21416 133912 117320 133940
rect 21416 133900 21422 133912
rect 117314 133900 117320 133912
rect 117372 133900 117378 133952
rect 14458 133832 14464 133884
rect 14516 133872 14522 133884
rect 117406 133872 117412 133884
rect 14516 133844 117412 133872
rect 14516 133832 14522 133844
rect 117406 133832 117412 133844
rect 117464 133832 117470 133884
rect 31018 132404 31024 132456
rect 31076 132444 31082 132456
rect 117314 132444 117320 132456
rect 31076 132416 117320 132444
rect 31076 132404 31082 132416
rect 117314 132404 117320 132416
rect 117372 132404 117378 132456
rect 18598 131044 18604 131096
rect 18656 131084 18662 131096
rect 117314 131084 117320 131096
rect 18656 131056 117320 131084
rect 18656 131044 18662 131056
rect 117314 131044 117320 131056
rect 117372 131044 117378 131096
rect 189166 129752 189172 129804
rect 189224 129792 189230 129804
rect 189626 129792 189632 129804
rect 189224 129764 189632 129792
rect 189224 129752 189230 129764
rect 189626 129752 189632 129764
rect 189684 129752 189690 129804
rect 13078 129684 13084 129736
rect 13136 129724 13142 129736
rect 117314 129724 117320 129736
rect 13136 129696 117320 129724
rect 13136 129684 13142 129696
rect 117314 129684 117320 129696
rect 117372 129684 117378 129736
rect 84930 128256 84936 128308
rect 84988 128296 84994 128308
rect 117314 128296 117320 128308
rect 84988 128268 117320 128296
rect 84988 128256 84994 128268
rect 117314 128256 117320 128268
rect 117372 128256 117378 128308
rect 10318 126896 10324 126948
rect 10376 126936 10382 126948
rect 117314 126936 117320 126948
rect 10376 126908 117320 126936
rect 10376 126896 10382 126908
rect 117314 126896 117320 126908
rect 117372 126896 117378 126948
rect 189258 126896 189264 126948
rect 189316 126936 189322 126948
rect 189626 126936 189632 126948
rect 189316 126908 189632 126936
rect 189316 126896 189322 126908
rect 189626 126896 189632 126908
rect 189684 126896 189690 126948
rect 48958 124108 48964 124160
rect 49016 124148 49022 124160
rect 117314 124148 117320 124160
rect 49016 124120 117320 124148
rect 49016 124108 49022 124120
rect 117314 124108 117320 124120
rect 117372 124108 117378 124160
rect 8938 122748 8944 122800
rect 8996 122788 9002 122800
rect 117314 122788 117320 122800
rect 8996 122760 117320 122788
rect 8996 122748 9002 122760
rect 117314 122748 117320 122760
rect 117372 122748 117378 122800
rect 17218 121388 17224 121440
rect 17276 121428 17282 121440
rect 117314 121428 117320 121440
rect 17276 121400 117320 121428
rect 17276 121388 17282 121400
rect 117314 121388 117320 121400
rect 117372 121388 117378 121440
rect 189074 121388 189080 121440
rect 189132 121428 189138 121440
rect 189350 121428 189356 121440
rect 189132 121400 189356 121428
rect 189132 121388 189138 121400
rect 189350 121388 189356 121400
rect 189408 121388 189414 121440
rect 7558 120028 7564 120080
rect 7616 120068 7622 120080
rect 117314 120068 117320 120080
rect 7616 120040 117320 120068
rect 7616 120028 7622 120040
rect 117314 120028 117320 120040
rect 117372 120028 117378 120080
rect 4798 118600 4804 118652
rect 4856 118640 4862 118652
rect 117314 118640 117320 118652
rect 4856 118612 117320 118640
rect 4856 118600 4862 118612
rect 117314 118600 117320 118612
rect 117372 118600 117378 118652
rect 40034 117240 40040 117292
rect 40092 117280 40098 117292
rect 117314 117280 117320 117292
rect 40092 117252 117320 117280
rect 40092 117240 40098 117252
rect 117314 117240 117320 117252
rect 117372 117240 117378 117292
rect 106918 115880 106924 115932
rect 106976 115920 106982 115932
rect 117314 115920 117320 115932
rect 106976 115892 117320 115920
rect 106976 115880 106982 115892
rect 117314 115880 117320 115892
rect 117372 115880 117378 115932
rect 189718 111800 189724 111852
rect 189776 111840 189782 111852
rect 580074 111840 580080 111852
rect 189776 111812 580080 111840
rect 189776 111800 189782 111812
rect 580074 111800 580080 111812
rect 580132 111800 580138 111852
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 21358 111772 21364 111784
rect 3384 111744 21364 111772
rect 3384 111732 3390 111744
rect 21358 111732 21364 111744
rect 21416 111732 21422 111784
rect 191926 108944 191932 108996
rect 191984 108984 191990 108996
rect 207658 108984 207664 108996
rect 191984 108956 207664 108984
rect 191984 108944 191990 108956
rect 207658 108944 207664 108956
rect 207716 108944 207722 108996
rect 191926 107584 191932 107636
rect 191984 107624 191990 107636
rect 206278 107624 206284 107636
rect 191984 107596 206284 107624
rect 191984 107584 191990 107596
rect 206278 107584 206284 107596
rect 206336 107584 206342 107636
rect 191926 106224 191932 106276
rect 191984 106264 191990 106276
rect 203518 106264 203524 106276
rect 191984 106236 203524 106264
rect 191984 106224 191990 106236
rect 203518 106224 203524 106236
rect 203576 106224 203582 106276
rect 193122 104796 193128 104848
rect 193180 104836 193186 104848
rect 200758 104836 200764 104848
rect 193180 104808 200764 104836
rect 193180 104796 193186 104808
rect 200758 104796 200764 104808
rect 200816 104796 200822 104848
rect 193122 102484 193128 102536
rect 193180 102524 193186 102536
rect 199378 102524 199384 102536
rect 193180 102496 199384 102524
rect 193180 102484 193186 102496
rect 199378 102484 199384 102496
rect 199436 102484 199442 102536
rect 191926 101124 191932 101176
rect 191984 101164 191990 101176
rect 197998 101164 198004 101176
rect 191984 101136 198004 101164
rect 191984 101124 191990 101136
rect 197998 101124 198004 101136
rect 198056 101124 198062 101176
rect 192386 100648 192392 100700
rect 192444 100688 192450 100700
rect 196618 100688 196624 100700
rect 192444 100660 196624 100688
rect 192444 100648 192450 100660
rect 196618 100648 196624 100660
rect 196676 100648 196682 100700
rect 192110 98472 192116 98524
rect 192168 98512 192174 98524
rect 193950 98512 193956 98524
rect 192168 98484 193956 98512
rect 192168 98472 192174 98484
rect 193950 98472 193956 98484
rect 194008 98472 194014 98524
rect 192202 97452 192208 97504
rect 192260 97492 192266 97504
rect 194042 97492 194048 97504
rect 192260 97464 194048 97492
rect 192260 97452 192266 97464
rect 194042 97452 194048 97464
rect 194100 97452 194106 97504
rect 191926 96432 191932 96484
rect 191984 96472 191990 96484
rect 194134 96472 194140 96484
rect 191984 96444 194140 96472
rect 191984 96432 191990 96444
rect 194134 96432 194140 96444
rect 194192 96432 194198 96484
rect 193122 95140 193128 95192
rect 193180 95180 193186 95192
rect 221458 95180 221464 95192
rect 193180 95152 221464 95180
rect 193180 95140 193186 95152
rect 221458 95140 221464 95152
rect 221516 95140 221522 95192
rect 360930 94528 360936 94580
rect 360988 94568 360994 94580
rect 580166 94568 580172 94580
rect 360988 94540 580172 94568
rect 360988 94528 360994 94540
rect 580166 94528 580172 94540
rect 580224 94528 580230 94580
rect 359550 94460 359556 94512
rect 359608 94500 359614 94512
rect 579982 94500 579988 94512
rect 359608 94472 579988 94500
rect 359608 94460 359614 94472
rect 579982 94460 579988 94472
rect 580040 94460 580046 94512
rect 193122 92420 193128 92472
rect 193180 92460 193186 92472
rect 360838 92460 360844 92472
rect 193180 92432 360844 92460
rect 193180 92420 193186 92432
rect 360838 92420 360844 92432
rect 360896 92420 360902 92472
rect 193122 90992 193128 91044
rect 193180 91032 193186 91044
rect 359458 91032 359464 91044
rect 193180 91004 359464 91032
rect 193180 90992 193186 91004
rect 359458 90992 359464 91004
rect 359516 90992 359522 91044
rect 193122 89632 193128 89684
rect 193180 89672 193186 89684
rect 202138 89672 202144 89684
rect 193180 89644 202144 89672
rect 193180 89632 193186 89644
rect 202138 89632 202144 89644
rect 202196 89632 202202 89684
rect 192938 88952 192944 89004
rect 192996 88992 193002 89004
rect 225598 88992 225604 89004
rect 192996 88964 225604 88992
rect 192996 88952 193002 88964
rect 225598 88952 225604 88964
rect 225656 88952 225662 89004
rect 193030 87592 193036 87644
rect 193088 87632 193094 87644
rect 224218 87632 224224 87644
rect 193088 87604 224224 87632
rect 193088 87592 193094 87604
rect 224218 87592 224224 87604
rect 224276 87592 224282 87644
rect 580166 86368 580172 86420
rect 580224 86408 580230 86420
rect 580810 86408 580816 86420
rect 580224 86380 580816 86408
rect 580224 86368 580230 86380
rect 580810 86368 580816 86380
rect 580868 86368 580874 86420
rect 193122 85484 193128 85536
rect 193180 85524 193186 85536
rect 360930 85524 360936 85536
rect 193180 85496 360936 85524
rect 193180 85484 193186 85496
rect 360930 85484 360936 85496
rect 360988 85484 360994 85536
rect 3326 84192 3332 84244
rect 3384 84232 3390 84244
rect 120626 84232 120632 84244
rect 3384 84204 120632 84232
rect 3384 84192 3390 84204
rect 120626 84192 120632 84204
rect 120684 84192 120690 84244
rect 193122 84124 193128 84176
rect 193180 84164 193186 84176
rect 359550 84164 359556 84176
rect 193180 84136 359556 84164
rect 193180 84124 193186 84136
rect 359550 84124 359556 84136
rect 359608 84124 359614 84176
rect 189074 80724 189080 80776
rect 189132 80764 189138 80776
rect 580258 80764 580264 80776
rect 189132 80736 580264 80764
rect 189132 80724 189138 80736
rect 580258 80724 580264 80736
rect 580316 80724 580322 80776
rect 188982 80656 188988 80708
rect 189040 80696 189046 80708
rect 580350 80696 580356 80708
rect 189040 80668 580356 80696
rect 189040 80656 189046 80668
rect 580350 80656 580356 80668
rect 580408 80656 580414 80708
rect 193122 80112 193128 80164
rect 193180 80152 193186 80164
rect 526438 80152 526444 80164
rect 193180 80124 526444 80152
rect 193180 80112 193186 80124
rect 526438 80112 526444 80124
rect 526496 80112 526502 80164
rect 127176 80056 131160 80084
rect 3694 79976 3700 80028
rect 3752 80016 3758 80028
rect 127066 80016 127072 80028
rect 3752 79988 127072 80016
rect 3752 79976 3758 79988
rect 127066 79976 127072 79988
rect 127124 79976 127130 80028
rect 127176 79960 127204 80056
rect 127250 79976 127256 80028
rect 127308 80016 127314 80028
rect 130194 80016 130200 80028
rect 127308 79988 130200 80016
rect 127308 79976 127314 79988
rect 130194 79976 130200 79988
rect 130252 79976 130258 80028
rect 131132 80016 131160 80056
rect 132926 80056 142982 80084
rect 131132 79988 131574 80016
rect 131546 79960 131574 79988
rect 131638 79988 132862 80016
rect 127158 79908 127164 79960
rect 127216 79908 127222 79960
rect 129918 79908 129924 79960
rect 129976 79948 129982 79960
rect 130792 79948 130798 79960
rect 129976 79920 130798 79948
rect 129976 79908 129982 79920
rect 130792 79908 130798 79920
rect 130850 79908 130856 79960
rect 130976 79908 130982 79960
rect 131034 79908 131040 79960
rect 131528 79908 131534 79960
rect 131586 79908 131592 79960
rect 121086 79840 121092 79892
rect 121144 79880 121150 79892
rect 129458 79880 129464 79892
rect 121144 79852 129464 79880
rect 121144 79840 121150 79852
rect 129458 79840 129464 79852
rect 129516 79840 129522 79892
rect 129550 79840 129556 79892
rect 129608 79880 129614 79892
rect 130994 79880 131022 79908
rect 129608 79852 131022 79880
rect 129608 79840 129614 79852
rect 131252 79840 131258 79892
rect 131310 79840 131316 79892
rect 126882 79772 126888 79824
rect 126940 79812 126946 79824
rect 131160 79812 131166 79824
rect 126940 79784 131166 79812
rect 126940 79772 126946 79784
rect 131160 79772 131166 79784
rect 131218 79772 131224 79824
rect 131022 79704 131028 79756
rect 131080 79744 131086 79756
rect 131270 79744 131298 79840
rect 131344 79772 131350 79824
rect 131402 79772 131408 79824
rect 131080 79716 131298 79744
rect 131080 79704 131086 79716
rect 126330 79636 126336 79688
rect 126388 79676 126394 79688
rect 126388 79648 127756 79676
rect 126388 79636 126394 79648
rect 119430 79568 119436 79620
rect 119488 79608 119494 79620
rect 127618 79608 127624 79620
rect 119488 79580 127624 79608
rect 119488 79568 119494 79580
rect 127618 79568 127624 79580
rect 127676 79568 127682 79620
rect 127728 79608 127756 79648
rect 131114 79636 131120 79688
rect 131172 79676 131178 79688
rect 131362 79676 131390 79772
rect 131172 79648 131390 79676
rect 131172 79636 131178 79648
rect 131638 79608 131666 79988
rect 131988 79908 131994 79960
rect 132046 79908 132052 79960
rect 131712 79840 131718 79892
rect 131770 79840 131776 79892
rect 131896 79840 131902 79892
rect 131954 79840 131960 79892
rect 131730 79676 131758 79840
rect 131914 79756 131942 79840
rect 131850 79704 131856 79756
rect 131908 79716 131942 79756
rect 132006 79744 132034 79908
rect 132834 79892 132862 79988
rect 132264 79840 132270 79892
rect 132322 79880 132328 79892
rect 132322 79852 132448 79880
rect 132322 79840 132328 79852
rect 132420 79812 132448 79852
rect 132816 79840 132822 79892
rect 132874 79840 132880 79892
rect 132374 79784 132448 79812
rect 132006 79716 132264 79744
rect 131908 79704 131914 79716
rect 131942 79676 131948 79688
rect 131730 79648 131948 79676
rect 131942 79636 131948 79648
rect 132000 79636 132006 79688
rect 132236 79620 132264 79716
rect 127728 79580 131666 79608
rect 132218 79568 132224 79620
rect 132276 79568 132282 79620
rect 132374 79608 132402 79784
rect 132540 79772 132546 79824
rect 132598 79812 132604 79824
rect 132926 79812 132954 80056
rect 142954 80016 142982 80056
rect 143138 80056 149146 80084
rect 143138 80016 143166 80056
rect 149118 80016 149146 80056
rect 149210 80056 149790 80084
rect 149210 80016 149238 80056
rect 136330 79988 140912 80016
rect 133368 79908 133374 79960
rect 133426 79908 133432 79960
rect 133552 79908 133558 79960
rect 133610 79908 133616 79960
rect 133736 79908 133742 79960
rect 133794 79908 133800 79960
rect 133828 79908 133834 79960
rect 133886 79908 133892 79960
rect 134196 79948 134202 79960
rect 133984 79920 134202 79948
rect 133184 79880 133190 79892
rect 132598 79772 132632 79812
rect 132604 79688 132632 79772
rect 132696 79784 132954 79812
rect 133018 79852 133190 79880
rect 132696 79688 132724 79784
rect 133018 79744 133046 79852
rect 133184 79840 133190 79852
rect 133242 79840 133248 79892
rect 132880 79716 133046 79744
rect 132880 79688 132908 79716
rect 133386 79688 133414 79908
rect 133570 79812 133598 79908
rect 133754 79824 133782 79908
rect 133524 79784 133598 79812
rect 133524 79756 133552 79784
rect 133690 79772 133696 79824
rect 133748 79784 133782 79824
rect 133748 79772 133754 79784
rect 133506 79704 133512 79756
rect 133564 79704 133570 79756
rect 133846 79688 133874 79908
rect 132586 79636 132592 79688
rect 132644 79636 132650 79688
rect 132678 79636 132684 79688
rect 132736 79636 132742 79688
rect 132862 79636 132868 79688
rect 132920 79636 132926 79688
rect 133322 79636 133328 79688
rect 133380 79648 133414 79688
rect 133380 79636 133386 79648
rect 133782 79636 133788 79688
rect 133840 79648 133874 79688
rect 133840 79636 133846 79648
rect 132494 79608 132500 79620
rect 132374 79580 132500 79608
rect 132494 79568 132500 79580
rect 132552 79568 132558 79620
rect 133984 79608 134012 79920
rect 134196 79908 134202 79920
rect 134254 79908 134260 79960
rect 135208 79908 135214 79960
rect 135266 79908 135272 79960
rect 134656 79840 134662 79892
rect 134714 79840 134720 79892
rect 134932 79840 134938 79892
rect 134990 79840 134996 79892
rect 135116 79840 135122 79892
rect 135174 79840 135180 79892
rect 134058 79636 134064 79688
rect 134116 79676 134122 79688
rect 134674 79676 134702 79840
rect 134116 79648 134702 79676
rect 134116 79636 134122 79648
rect 134794 79636 134800 79688
rect 134852 79676 134858 79688
rect 134950 79676 134978 79840
rect 135134 79744 135162 79840
rect 135088 79716 135162 79744
rect 135088 79688 135116 79716
rect 135226 79688 135254 79908
rect 135852 79880 135858 79892
rect 135732 79852 135858 79880
rect 134852 79648 134978 79676
rect 134852 79636 134858 79648
rect 135070 79636 135076 79688
rect 135128 79636 135134 79688
rect 135162 79636 135168 79688
rect 135220 79648 135254 79688
rect 135220 79636 135226 79648
rect 135622 79636 135628 79688
rect 135680 79676 135686 79688
rect 135732 79676 135760 79852
rect 135852 79840 135858 79852
rect 135910 79840 135916 79892
rect 135944 79840 135950 79892
rect 136002 79840 136008 79892
rect 135680 79648 135760 79676
rect 135962 79676 135990 79840
rect 135962 79648 136036 79676
rect 135680 79636 135686 79648
rect 134150 79608 134156 79620
rect 133984 79580 134156 79608
rect 134150 79568 134156 79580
rect 134208 79568 134214 79620
rect 135898 79608 135904 79620
rect 135226 79580 135904 79608
rect 120626 79500 120632 79552
rect 120684 79540 120690 79552
rect 129366 79540 129372 79552
rect 120684 79512 129372 79540
rect 120684 79500 120690 79512
rect 129366 79500 129372 79512
rect 129424 79500 129430 79552
rect 129458 79500 129464 79552
rect 129516 79540 129522 79552
rect 135226 79540 135254 79580
rect 135898 79568 135904 79580
rect 135956 79568 135962 79620
rect 129516 79512 135254 79540
rect 129516 79500 129522 79512
rect 135438 79500 135444 79552
rect 135496 79540 135502 79552
rect 136008 79540 136036 79648
rect 135496 79512 136036 79540
rect 135496 79500 135502 79512
rect 136330 79484 136358 79988
rect 136680 79908 136686 79960
rect 136738 79908 136744 79960
rect 136772 79908 136778 79960
rect 136830 79908 136836 79960
rect 136864 79908 136870 79960
rect 136922 79948 136928 79960
rect 136922 79908 136956 79948
rect 137508 79908 137514 79960
rect 137566 79908 137572 79960
rect 138152 79908 138158 79960
rect 138210 79908 138216 79960
rect 139532 79948 139538 79960
rect 138308 79920 139118 79948
rect 136588 79880 136594 79892
rect 136560 79840 136594 79880
rect 136646 79840 136652 79892
rect 136560 79688 136588 79840
rect 136698 79756 136726 79908
rect 136790 79880 136818 79908
rect 136790 79852 136864 79880
rect 136836 79824 136864 79852
rect 136818 79772 136824 79824
rect 136876 79772 136882 79824
rect 136698 79716 136732 79756
rect 136726 79704 136732 79716
rect 136784 79704 136790 79756
rect 136542 79636 136548 79688
rect 136600 79636 136606 79688
rect 116670 79432 116676 79484
rect 116728 79472 116734 79484
rect 116728 79444 118694 79472
rect 116728 79432 116734 79444
rect 118666 79404 118694 79444
rect 127618 79432 127624 79484
rect 127676 79472 127682 79484
rect 135346 79472 135352 79484
rect 127676 79444 135352 79472
rect 127676 79432 127682 79444
rect 135346 79432 135352 79444
rect 135404 79432 135410 79484
rect 136266 79432 136272 79484
rect 136324 79444 136358 79484
rect 136928 79472 136956 79908
rect 137526 79744 137554 79908
rect 137876 79840 137882 79892
rect 137934 79840 137940 79892
rect 137020 79716 137554 79744
rect 137020 79552 137048 79716
rect 137094 79636 137100 79688
rect 137152 79676 137158 79688
rect 137894 79676 137922 79840
rect 137152 79648 137922 79676
rect 137152 79636 137158 79648
rect 138014 79636 138020 79688
rect 138072 79676 138078 79688
rect 138170 79676 138198 79908
rect 138308 79688 138336 79920
rect 139090 79892 139118 79920
rect 139182 79920 139538 79948
rect 138888 79880 138894 79892
rect 138492 79852 138894 79880
rect 138492 79688 138520 79852
rect 138888 79840 138894 79852
rect 138946 79840 138952 79892
rect 139072 79840 139078 79892
rect 139130 79840 139136 79892
rect 139182 79688 139210 79920
rect 139532 79908 139538 79920
rect 139590 79908 139596 79960
rect 140360 79948 140366 79960
rect 139918 79920 140366 79948
rect 139256 79840 139262 79892
rect 139314 79840 139320 79892
rect 139716 79880 139722 79892
rect 139596 79852 139722 79880
rect 138072 79648 138198 79676
rect 138072 79636 138078 79648
rect 138290 79636 138296 79688
rect 138348 79636 138354 79688
rect 138474 79636 138480 79688
rect 138532 79636 138538 79688
rect 139118 79636 139124 79688
rect 139176 79648 139210 79688
rect 139176 79636 139182 79648
rect 139274 79620 139302 79840
rect 139596 79688 139624 79852
rect 139716 79840 139722 79852
rect 139774 79840 139780 79892
rect 139808 79812 139814 79824
rect 139688 79784 139814 79812
rect 139578 79636 139584 79688
rect 139636 79636 139642 79688
rect 139210 79568 139216 79620
rect 139268 79580 139302 79620
rect 139688 79608 139716 79784
rect 139808 79772 139814 79784
rect 139866 79772 139872 79824
rect 139412 79580 139716 79608
rect 139268 79568 139274 79580
rect 139412 79552 139440 79580
rect 137002 79500 137008 79552
rect 137060 79500 137066 79552
rect 139394 79500 139400 79552
rect 139452 79500 139458 79552
rect 137738 79472 137744 79484
rect 136928 79444 137744 79472
rect 136324 79432 136330 79444
rect 137738 79432 137744 79444
rect 137796 79432 137802 79484
rect 139762 79432 139768 79484
rect 139820 79472 139826 79484
rect 139918 79472 139946 79920
rect 140360 79908 140366 79920
rect 140418 79908 140424 79960
rect 140452 79908 140458 79960
rect 140510 79908 140516 79960
rect 140544 79908 140550 79960
rect 140602 79908 140608 79960
rect 140084 79840 140090 79892
rect 140142 79840 140148 79892
rect 140176 79840 140182 79892
rect 140234 79840 140240 79892
rect 140102 79620 140130 79840
rect 140194 79688 140222 79840
rect 140314 79772 140320 79824
rect 140372 79812 140378 79824
rect 140470 79812 140498 79908
rect 140372 79784 140498 79812
rect 140372 79772 140378 79784
rect 140406 79704 140412 79756
rect 140464 79744 140470 79756
rect 140562 79744 140590 79908
rect 140636 79840 140642 79892
rect 140694 79840 140700 79892
rect 140884 79880 140912 79988
rect 141160 79988 141510 80016
rect 141004 79880 141010 79892
rect 140884 79852 141010 79880
rect 141004 79840 141010 79852
rect 141062 79840 141068 79892
rect 140464 79716 140590 79744
rect 140464 79704 140470 79716
rect 140194 79648 140228 79688
rect 140222 79636 140228 79648
rect 140280 79636 140286 79688
rect 140038 79568 140044 79620
rect 140096 79580 140130 79620
rect 140654 79608 140682 79840
rect 141160 79620 141188 79988
rect 141482 79960 141510 79988
rect 141620 79988 142062 80016
rect 142954 79988 143166 80016
rect 143782 79988 144086 80016
rect 141372 79948 141378 79960
rect 141252 79920 141378 79948
rect 141252 79688 141280 79920
rect 141372 79908 141378 79920
rect 141430 79908 141436 79960
rect 141464 79908 141470 79960
rect 141522 79908 141528 79960
rect 141234 79636 141240 79688
rect 141292 79636 141298 79688
rect 140774 79608 140780 79620
rect 140424 79580 140682 79608
rect 140096 79568 140102 79580
rect 139820 79444 139946 79472
rect 140424 79472 140452 79580
rect 140746 79568 140780 79608
rect 140832 79568 140838 79620
rect 141142 79568 141148 79620
rect 141200 79568 141206 79620
rect 140498 79500 140504 79552
rect 140556 79540 140562 79552
rect 140746 79540 140774 79568
rect 140556 79512 140774 79540
rect 140556 79500 140562 79512
rect 141050 79500 141056 79552
rect 141108 79540 141114 79552
rect 141620 79540 141648 79988
rect 142034 79960 142062 79988
rect 143782 79960 143810 79988
rect 141740 79908 141746 79960
rect 141798 79908 141804 79960
rect 141832 79908 141838 79960
rect 141890 79908 141896 79960
rect 141924 79908 141930 79960
rect 141982 79908 141988 79960
rect 142016 79908 142022 79960
rect 142074 79908 142080 79960
rect 142108 79908 142114 79960
rect 142166 79908 142172 79960
rect 142292 79948 142298 79960
rect 142264 79908 142298 79948
rect 142350 79908 142356 79960
rect 142752 79908 142758 79960
rect 142810 79908 142816 79960
rect 142936 79908 142942 79960
rect 142994 79908 143000 79960
rect 143028 79908 143034 79960
rect 143086 79948 143092 79960
rect 143086 79920 143718 79948
rect 143086 79908 143092 79920
rect 141758 79824 141786 79908
rect 141694 79772 141700 79824
rect 141752 79784 141786 79824
rect 141752 79772 141758 79784
rect 141850 79688 141878 79908
rect 141942 79744 141970 79908
rect 141942 79716 142016 79744
rect 141850 79648 141884 79688
rect 141878 79636 141884 79648
rect 141936 79636 141942 79688
rect 141108 79512 141648 79540
rect 141108 79500 141114 79512
rect 140774 79472 140780 79484
rect 140424 79444 140780 79472
rect 139820 79432 139826 79444
rect 140774 79432 140780 79444
rect 140832 79432 140838 79484
rect 141786 79432 141792 79484
rect 141844 79472 141850 79484
rect 141988 79472 142016 79716
rect 142126 79688 142154 79908
rect 142264 79688 142292 79908
rect 142384 79880 142390 79892
rect 142356 79840 142390 79880
rect 142442 79840 142448 79892
rect 142476 79840 142482 79892
rect 142534 79840 142540 79892
rect 142568 79840 142574 79892
rect 142626 79840 142632 79892
rect 142356 79756 142384 79840
rect 142338 79704 142344 79756
rect 142396 79704 142402 79756
rect 142062 79636 142068 79688
rect 142120 79648 142154 79688
rect 142120 79636 142126 79648
rect 142246 79636 142252 79688
rect 142304 79636 142310 79688
rect 142494 79608 142522 79840
rect 142586 79676 142614 79840
rect 142770 79744 142798 79908
rect 142954 79824 142982 79908
rect 143580 79840 143586 79892
rect 143638 79840 143644 79892
rect 142954 79784 142988 79824
rect 142982 79772 142988 79784
rect 143040 79772 143046 79824
rect 143598 79756 143626 79840
rect 143690 79824 143718 79920
rect 143764 79908 143770 79960
rect 143822 79908 143828 79960
rect 143948 79880 143954 79892
rect 143828 79852 143954 79880
rect 143690 79784 143724 79824
rect 143718 79772 143724 79784
rect 143776 79772 143782 79824
rect 142770 79716 143488 79744
rect 143598 79716 143632 79756
rect 143460 79688 143488 79716
rect 143626 79704 143632 79716
rect 143684 79704 143690 79756
rect 142706 79676 142712 79688
rect 142586 79648 142712 79676
rect 142706 79636 142712 79648
rect 142764 79636 142770 79688
rect 142890 79636 142896 79688
rect 142948 79636 142954 79688
rect 143442 79636 143448 79688
rect 143500 79636 143506 79688
rect 143534 79636 143540 79688
rect 143592 79676 143598 79688
rect 143828 79676 143856 79852
rect 143948 79840 143954 79852
rect 144006 79840 144012 79892
rect 144058 79744 144086 79988
rect 144978 79988 147214 80016
rect 149118 79988 149238 80016
rect 149762 80016 149790 80056
rect 149900 80056 170490 80084
rect 149900 80016 149928 80056
rect 170462 80016 170490 80056
rect 172486 80056 174906 80084
rect 172486 80016 172514 80056
rect 174878 80016 174906 80056
rect 175062 80056 178494 80084
rect 175062 80016 175090 80056
rect 149762 79988 149928 80016
rect 153764 79988 154206 80016
rect 144776 79948 144782 79960
rect 143592 79648 143856 79676
rect 143966 79716 144086 79744
rect 144150 79920 144782 79948
rect 143592 79636 143598 79648
rect 141844 79444 142016 79472
rect 142356 79580 142522 79608
rect 142356 79472 142384 79580
rect 142430 79500 142436 79552
rect 142488 79540 142494 79552
rect 142908 79540 142936 79636
rect 143966 79620 143994 79716
rect 144150 79676 144178 79920
rect 144776 79908 144782 79920
rect 144834 79908 144840 79960
rect 144868 79908 144874 79960
rect 144926 79908 144932 79960
rect 144408 79840 144414 79892
rect 144466 79840 144472 79892
rect 144500 79840 144506 79892
rect 144558 79880 144564 79892
rect 144558 79852 144776 79880
rect 144558 79840 144564 79852
rect 143902 79568 143908 79620
rect 143960 79580 143994 79620
rect 144104 79648 144178 79676
rect 143960 79568 143966 79580
rect 144104 79552 144132 79648
rect 144426 79608 144454 79840
rect 144748 79824 144776 79852
rect 144886 79824 144914 79908
rect 144730 79772 144736 79824
rect 144788 79772 144794 79824
rect 144822 79772 144828 79824
rect 144880 79784 144914 79824
rect 144880 79772 144886 79784
rect 144638 79608 144644 79620
rect 144426 79580 144644 79608
rect 144638 79568 144644 79580
rect 144696 79568 144702 79620
rect 142488 79512 142936 79540
rect 142488 79500 142494 79512
rect 144086 79500 144092 79552
rect 144144 79500 144150 79552
rect 142890 79472 142896 79484
rect 142356 79444 142896 79472
rect 141844 79432 141850 79444
rect 142890 79432 142896 79444
rect 142948 79432 142954 79484
rect 144362 79432 144368 79484
rect 144420 79472 144426 79484
rect 144978 79472 145006 79988
rect 147186 79960 147214 79988
rect 145236 79908 145242 79960
rect 145294 79908 145300 79960
rect 145512 79908 145518 79960
rect 145570 79908 145576 79960
rect 146984 79948 146990 79960
rect 146542 79920 146990 79948
rect 145052 79772 145058 79824
rect 145110 79772 145116 79824
rect 144420 79444 145006 79472
rect 145070 79472 145098 79772
rect 145254 79552 145282 79908
rect 145254 79512 145288 79552
rect 145282 79500 145288 79512
rect 145340 79500 145346 79552
rect 145190 79472 145196 79484
rect 145070 79444 145196 79472
rect 144420 79432 144426 79444
rect 145190 79432 145196 79444
rect 145248 79432 145254 79484
rect 145530 79472 145558 79908
rect 146156 79840 146162 79892
rect 146214 79840 146220 79892
rect 146248 79840 146254 79892
rect 146306 79840 146312 79892
rect 146340 79840 146346 79892
rect 146398 79840 146404 79892
rect 146174 79688 146202 79840
rect 146266 79744 146294 79840
rect 146358 79812 146386 79840
rect 146358 79784 146432 79812
rect 146266 79716 146340 79744
rect 146174 79648 146208 79688
rect 146202 79636 146208 79648
rect 146260 79636 146266 79688
rect 145650 79500 145656 79552
rect 145708 79540 145714 79552
rect 146312 79540 146340 79716
rect 145708 79512 146340 79540
rect 146404 79540 146432 79784
rect 146542 79744 146570 79920
rect 146984 79908 146990 79920
rect 147042 79908 147048 79960
rect 147168 79908 147174 79960
rect 147226 79908 147232 79960
rect 147904 79948 147910 79960
rect 147646 79920 147910 79948
rect 146616 79840 146622 79892
rect 146674 79840 146680 79892
rect 146800 79840 146806 79892
rect 146858 79880 146864 79892
rect 146858 79852 147076 79880
rect 146858 79840 146864 79852
rect 146634 79812 146662 79840
rect 146634 79784 146984 79812
rect 146542 79716 146892 79744
rect 146754 79540 146760 79552
rect 146404 79512 146760 79540
rect 145708 79500 145714 79512
rect 146754 79500 146760 79512
rect 146812 79500 146818 79552
rect 145926 79472 145932 79484
rect 145530 79444 145932 79472
rect 145926 79432 145932 79444
rect 145984 79432 145990 79484
rect 146294 79432 146300 79484
rect 146352 79472 146358 79484
rect 146864 79472 146892 79716
rect 146956 79688 146984 79784
rect 146938 79636 146944 79688
rect 146996 79636 147002 79688
rect 146352 79444 146892 79472
rect 146352 79432 146358 79444
rect 144914 79404 144920 79416
rect 118666 79376 144920 79404
rect 144914 79364 144920 79376
rect 144972 79364 144978 79416
rect 145098 79364 145104 79416
rect 145156 79404 145162 79416
rect 145834 79404 145840 79416
rect 145156 79376 145840 79404
rect 145156 79364 145162 79376
rect 145834 79364 145840 79376
rect 145892 79364 145898 79416
rect 146478 79364 146484 79416
rect 146536 79404 146542 79416
rect 147048 79404 147076 79852
rect 147260 79840 147266 79892
rect 147318 79840 147324 79892
rect 147352 79840 147358 79892
rect 147410 79880 147416 79892
rect 147410 79840 147444 79880
rect 147278 79688 147306 79840
rect 147416 79756 147444 79840
rect 147536 79772 147542 79824
rect 147594 79772 147600 79824
rect 147398 79704 147404 79756
rect 147456 79704 147462 79756
rect 147554 79688 147582 79772
rect 147214 79636 147220 79688
rect 147272 79648 147306 79688
rect 147272 79636 147278 79648
rect 147490 79636 147496 79688
rect 147548 79648 147582 79688
rect 147548 79636 147554 79648
rect 147122 79568 147128 79620
rect 147180 79608 147186 79620
rect 147646 79608 147674 79920
rect 147904 79908 147910 79920
rect 147962 79908 147968 79960
rect 148180 79908 148186 79960
rect 148238 79908 148244 79960
rect 148272 79908 148278 79960
rect 148330 79908 148336 79960
rect 148364 79908 148370 79960
rect 148422 79908 148428 79960
rect 148732 79948 148738 79960
rect 148704 79908 148738 79948
rect 148790 79908 148796 79960
rect 149376 79908 149382 79960
rect 149434 79948 149440 79960
rect 149434 79908 149468 79948
rect 149928 79908 149934 79960
rect 149986 79908 149992 79960
rect 150020 79908 150026 79960
rect 150078 79908 150084 79960
rect 151124 79948 151130 79960
rect 150912 79920 151130 79948
rect 147812 79840 147818 79892
rect 147870 79880 147876 79892
rect 147870 79852 147950 79880
rect 147870 79840 147876 79852
rect 147720 79772 147726 79824
rect 147778 79772 147784 79824
rect 147738 79688 147766 79772
rect 147738 79648 147772 79688
rect 147766 79636 147772 79648
rect 147824 79636 147830 79688
rect 147180 79580 147674 79608
rect 147180 79568 147186 79580
rect 146536 79376 147076 79404
rect 147922 79404 147950 79852
rect 148198 79688 148226 79908
rect 148290 79756 148318 79908
rect 148382 79812 148410 79908
rect 148548 79840 148554 79892
rect 148606 79840 148612 79892
rect 148382 79784 148456 79812
rect 148290 79716 148324 79756
rect 148318 79704 148324 79716
rect 148376 79704 148382 79756
rect 148428 79688 148456 79784
rect 148198 79648 148232 79688
rect 148226 79636 148232 79648
rect 148284 79636 148290 79688
rect 148410 79636 148416 79688
rect 148468 79636 148474 79688
rect 148566 79620 148594 79840
rect 148704 79620 148732 79908
rect 148916 79880 148922 79892
rect 148796 79852 148922 79880
rect 148796 79824 148824 79852
rect 148916 79840 148922 79852
rect 148974 79840 148980 79892
rect 149008 79840 149014 79892
rect 149066 79840 149072 79892
rect 149192 79880 149198 79892
rect 149164 79840 149198 79880
rect 149250 79840 149256 79892
rect 149440 79880 149468 79908
rect 149440 79852 149560 79880
rect 148778 79772 148784 79824
rect 148836 79772 148842 79824
rect 148870 79704 148876 79756
rect 148928 79744 148934 79756
rect 149026 79744 149054 79840
rect 149164 79756 149192 79840
rect 148928 79716 149054 79744
rect 148928 79704 148934 79716
rect 149146 79704 149152 79756
rect 149204 79704 149210 79756
rect 149422 79636 149428 79688
rect 149480 79676 149486 79688
rect 149532 79676 149560 79852
rect 149652 79840 149658 79892
rect 149710 79840 149716 79892
rect 149480 79648 149560 79676
rect 149480 79636 149486 79648
rect 148566 79580 148600 79620
rect 148594 79568 148600 79580
rect 148652 79568 148658 79620
rect 148686 79568 148692 79620
rect 148744 79568 148750 79620
rect 149670 79540 149698 79840
rect 149946 79812 149974 79908
rect 149900 79784 149974 79812
rect 149900 79688 149928 79784
rect 150038 79756 150066 79908
rect 150204 79840 150210 79892
rect 150262 79840 150268 79892
rect 150388 79840 150394 79892
rect 150446 79840 150452 79892
rect 150480 79840 150486 79892
rect 150538 79840 150544 79892
rect 150664 79840 150670 79892
rect 150722 79880 150728 79892
rect 150722 79852 150848 79880
rect 150722 79840 150728 79852
rect 149974 79704 149980 79756
rect 150032 79716 150066 79756
rect 150032 79704 150038 79716
rect 150222 79688 150250 79840
rect 149882 79636 149888 79688
rect 149940 79636 149946 79688
rect 150222 79648 150256 79688
rect 150250 79636 150256 79648
rect 150308 79636 150314 79688
rect 150406 79608 150434 79840
rect 150498 79676 150526 79840
rect 150572 79772 150578 79824
rect 150630 79812 150636 79824
rect 150630 79784 150756 79812
rect 150630 79772 150636 79784
rect 150728 79756 150756 79784
rect 150710 79704 150716 79756
rect 150768 79704 150774 79756
rect 150618 79676 150624 79688
rect 150498 79648 150624 79676
rect 150618 79636 150624 79648
rect 150676 79636 150682 79688
rect 150360 79580 150434 79608
rect 150158 79540 150164 79552
rect 149670 79512 150164 79540
rect 150158 79500 150164 79512
rect 150216 79500 150222 79552
rect 149238 79432 149244 79484
rect 149296 79472 149302 79484
rect 149514 79472 149520 79484
rect 149296 79444 149520 79472
rect 149296 79432 149302 79444
rect 149514 79432 149520 79444
rect 149572 79432 149578 79484
rect 148962 79404 148968 79416
rect 147922 79376 148968 79404
rect 146536 79364 146542 79376
rect 148962 79364 148968 79376
rect 149020 79364 149026 79416
rect 149330 79364 149336 79416
rect 149388 79404 149394 79416
rect 149790 79404 149796 79416
rect 149388 79376 149796 79404
rect 149388 79364 149394 79376
rect 149790 79364 149796 79376
rect 149848 79364 149854 79416
rect 150360 79404 150388 79580
rect 150434 79500 150440 79552
rect 150492 79540 150498 79552
rect 150820 79540 150848 79852
rect 150912 79620 150940 79920
rect 151124 79908 151130 79920
rect 151182 79908 151188 79960
rect 151308 79908 151314 79960
rect 151366 79908 151372 79960
rect 151400 79908 151406 79960
rect 151458 79908 151464 79960
rect 151492 79908 151498 79960
rect 151550 79908 151556 79960
rect 151952 79908 151958 79960
rect 152010 79908 152016 79960
rect 152504 79908 152510 79960
rect 152562 79908 152568 79960
rect 152596 79908 152602 79960
rect 152654 79948 152660 79960
rect 152654 79908 152688 79948
rect 152780 79908 152786 79960
rect 152838 79908 152844 79960
rect 152964 79908 152970 79960
rect 153022 79908 153028 79960
rect 153056 79908 153062 79960
rect 153114 79908 153120 79960
rect 153148 79908 153154 79960
rect 153206 79908 153212 79960
rect 153240 79908 153246 79960
rect 153298 79908 153304 79960
rect 151032 79840 151038 79892
rect 151090 79880 151096 79892
rect 151216 79880 151222 79892
rect 151090 79840 151124 79880
rect 151096 79756 151124 79840
rect 151188 79840 151222 79880
rect 151274 79840 151280 79892
rect 151188 79756 151216 79840
rect 151326 79756 151354 79908
rect 151078 79704 151084 79756
rect 151136 79704 151142 79756
rect 151170 79704 151176 79756
rect 151228 79704 151234 79756
rect 151262 79704 151268 79756
rect 151320 79716 151354 79756
rect 151320 79704 151326 79716
rect 151418 79688 151446 79908
rect 151354 79636 151360 79688
rect 151412 79648 151446 79688
rect 151412 79636 151418 79648
rect 151510 79620 151538 79908
rect 151768 79840 151774 79892
rect 151826 79840 151832 79892
rect 151860 79840 151866 79892
rect 151918 79840 151924 79892
rect 151786 79812 151814 79840
rect 151648 79784 151814 79812
rect 151648 79620 151676 79784
rect 151878 79744 151906 79840
rect 151740 79716 151906 79744
rect 151740 79688 151768 79716
rect 151970 79688 151998 79908
rect 152228 79880 152234 79892
rect 151722 79636 151728 79688
rect 151780 79636 151786 79688
rect 151906 79636 151912 79688
rect 151964 79648 151998 79688
rect 152062 79852 152234 79880
rect 151964 79636 151970 79648
rect 150894 79568 150900 79620
rect 150952 79568 150958 79620
rect 151446 79568 151452 79620
rect 151504 79580 151538 79620
rect 151504 79568 151510 79580
rect 151630 79568 151636 79620
rect 151688 79568 151694 79620
rect 151814 79568 151820 79620
rect 151872 79608 151878 79620
rect 152062 79608 152090 79852
rect 152228 79840 152234 79852
rect 152286 79840 152292 79892
rect 152412 79880 152418 79892
rect 152384 79840 152418 79880
rect 152470 79840 152476 79892
rect 152136 79772 152142 79824
rect 152194 79812 152200 79824
rect 152194 79784 152320 79812
rect 152194 79772 152200 79784
rect 152292 79756 152320 79784
rect 152384 79756 152412 79840
rect 152274 79704 152280 79756
rect 152332 79704 152338 79756
rect 152366 79704 152372 79756
rect 152424 79704 152430 79756
rect 151872 79580 152090 79608
rect 152522 79620 152550 79908
rect 152660 79756 152688 79908
rect 152798 79756 152826 79908
rect 152642 79704 152648 79756
rect 152700 79704 152706 79756
rect 152798 79716 152832 79756
rect 152826 79704 152832 79716
rect 152884 79704 152890 79756
rect 152982 79676 153010 79908
rect 153074 79756 153102 79908
rect 153166 79812 153194 79908
rect 153258 79880 153286 79908
rect 153258 79852 153332 79880
rect 153166 79784 153240 79812
rect 153074 79716 153108 79756
rect 153102 79704 153108 79716
rect 153160 79704 153166 79756
rect 152660 79648 153010 79676
rect 152522 79580 152556 79620
rect 151872 79568 151878 79580
rect 152550 79568 152556 79580
rect 152608 79568 152614 79620
rect 150492 79512 150848 79540
rect 150492 79500 150498 79512
rect 152182 79500 152188 79552
rect 152240 79540 152246 79552
rect 152660 79540 152688 79648
rect 153212 79552 153240 79784
rect 153304 79688 153332 79852
rect 153516 79812 153522 79824
rect 153396 79784 153522 79812
rect 153286 79636 153292 79688
rect 153344 79636 153350 79688
rect 152240 79512 152688 79540
rect 152240 79500 152246 79512
rect 153194 79500 153200 79552
rect 153252 79500 153258 79552
rect 153010 79432 153016 79484
rect 153068 79472 153074 79484
rect 153396 79472 153424 79784
rect 153516 79772 153522 79784
rect 153574 79772 153580 79824
rect 153608 79772 153614 79824
rect 153666 79772 153672 79824
rect 153626 79688 153654 79772
rect 153562 79636 153568 79688
rect 153620 79648 153654 79688
rect 153620 79636 153626 79648
rect 153764 79552 153792 79988
rect 154178 79960 154206 79988
rect 156754 79988 157242 80016
rect 153884 79908 153890 79960
rect 153942 79908 153948 79960
rect 153976 79908 153982 79960
rect 154034 79908 154040 79960
rect 154068 79908 154074 79960
rect 154126 79908 154132 79960
rect 154160 79908 154166 79960
rect 154218 79908 154224 79960
rect 154252 79908 154258 79960
rect 154310 79908 154316 79960
rect 154344 79908 154350 79960
rect 154402 79948 154408 79960
rect 154402 79920 154482 79948
rect 154402 79908 154408 79920
rect 153902 79688 153930 79908
rect 153994 79756 154022 79908
rect 154086 79812 154114 79908
rect 154270 79880 154298 79908
rect 154270 79852 154344 79880
rect 154086 79784 154160 79812
rect 153994 79716 154028 79756
rect 154022 79704 154028 79716
rect 154080 79704 154086 79756
rect 153838 79636 153844 79688
rect 153896 79648 153930 79688
rect 153896 79636 153902 79648
rect 153930 79568 153936 79620
rect 153988 79608 153994 79620
rect 154132 79608 154160 79784
rect 154316 79756 154344 79852
rect 154454 79756 154482 79920
rect 154528 79908 154534 79960
rect 154586 79908 154592 79960
rect 154620 79908 154626 79960
rect 154678 79908 154684 79960
rect 154712 79908 154718 79960
rect 154770 79908 154776 79960
rect 154988 79908 154994 79960
rect 155046 79908 155052 79960
rect 155080 79908 155086 79960
rect 155138 79908 155144 79960
rect 155172 79908 155178 79960
rect 155230 79908 155236 79960
rect 155264 79908 155270 79960
rect 155322 79948 155328 79960
rect 155448 79948 155454 79960
rect 155322 79908 155356 79948
rect 154298 79704 154304 79756
rect 154356 79704 154362 79756
rect 154390 79704 154396 79756
rect 154448 79716 154482 79756
rect 154448 79704 154454 79716
rect 154546 79688 154574 79908
rect 154638 79756 154666 79908
rect 154730 79880 154758 79908
rect 154730 79852 154804 79880
rect 154638 79716 154672 79756
rect 154666 79704 154672 79716
rect 154724 79704 154730 79756
rect 154482 79636 154488 79688
rect 154540 79648 154574 79688
rect 154540 79636 154546 79648
rect 153988 79580 154160 79608
rect 153988 79568 153994 79580
rect 154574 79568 154580 79620
rect 154632 79608 154638 79620
rect 154776 79608 154804 79852
rect 155006 79756 155034 79908
rect 155098 79824 155126 79908
rect 155190 79880 155218 79908
rect 155190 79852 155264 79880
rect 155098 79784 155132 79824
rect 155126 79772 155132 79784
rect 155184 79772 155190 79824
rect 154942 79704 154948 79756
rect 155000 79716 155034 79756
rect 155000 79704 155006 79716
rect 154632 79580 154804 79608
rect 154632 79568 154638 79580
rect 155034 79568 155040 79620
rect 155092 79608 155098 79620
rect 155236 79608 155264 79852
rect 155092 79580 155264 79608
rect 155092 79568 155098 79580
rect 153746 79500 153752 79552
rect 153804 79500 153810 79552
rect 155218 79500 155224 79552
rect 155276 79540 155282 79552
rect 155328 79540 155356 79908
rect 155420 79908 155454 79948
rect 155506 79908 155512 79960
rect 155650 79920 155954 79948
rect 155420 79756 155448 79908
rect 155402 79704 155408 79756
rect 155460 79704 155466 79756
rect 155650 79688 155678 79920
rect 155926 79892 155954 79920
rect 156092 79908 156098 79960
rect 156150 79908 156156 79960
rect 156184 79908 156190 79960
rect 156242 79908 156248 79960
rect 156276 79908 156282 79960
rect 156334 79908 156340 79960
rect 155724 79840 155730 79892
rect 155782 79880 155788 79892
rect 155782 79840 155816 79880
rect 155908 79840 155914 79892
rect 155966 79840 155972 79892
rect 156000 79840 156006 79892
rect 156058 79840 156064 79892
rect 155650 79648 155684 79688
rect 155678 79636 155684 79648
rect 155736 79636 155742 79688
rect 155788 79552 155816 79840
rect 155862 79704 155868 79756
rect 155920 79744 155926 79756
rect 156018 79744 156046 79840
rect 155920 79716 156046 79744
rect 155920 79704 155926 79716
rect 156110 79620 156138 79908
rect 156202 79756 156230 79908
rect 156294 79812 156322 79908
rect 156368 79840 156374 79892
rect 156426 79880 156432 79892
rect 156552 79880 156558 79892
rect 156426 79840 156460 79880
rect 156294 79784 156368 79812
rect 156202 79716 156236 79756
rect 156230 79704 156236 79716
rect 156288 79704 156294 79756
rect 156340 79620 156368 79784
rect 156110 79580 156144 79620
rect 156138 79568 156144 79580
rect 156196 79568 156202 79620
rect 156322 79568 156328 79620
rect 156380 79568 156386 79620
rect 156432 79552 156460 79840
rect 156524 79840 156558 79880
rect 156610 79840 156616 79892
rect 156524 79620 156552 79840
rect 156754 79824 156782 79988
rect 157214 79960 157242 79988
rect 161722 79988 162440 80016
rect 161722 79960 161750 79988
rect 156828 79908 156834 79960
rect 156886 79908 156892 79960
rect 157104 79908 157110 79960
rect 157162 79908 157168 79960
rect 157196 79908 157202 79960
rect 157254 79908 157260 79960
rect 157380 79908 157386 79960
rect 157438 79908 157444 79960
rect 157472 79908 157478 79960
rect 157530 79908 157536 79960
rect 157564 79908 157570 79960
rect 157622 79908 157628 79960
rect 157656 79908 157662 79960
rect 157714 79948 157720 79960
rect 157714 79920 157978 79948
rect 157714 79908 157720 79920
rect 156846 79880 156874 79908
rect 156846 79852 156920 79880
rect 156754 79784 156788 79824
rect 156782 79772 156788 79784
rect 156840 79772 156846 79824
rect 156506 79568 156512 79620
rect 156564 79568 156570 79620
rect 155276 79512 155356 79540
rect 155276 79500 155282 79512
rect 155770 79500 155776 79552
rect 155828 79500 155834 79552
rect 156414 79500 156420 79552
rect 156472 79500 156478 79552
rect 156598 79500 156604 79552
rect 156656 79540 156662 79552
rect 156892 79540 156920 79852
rect 157122 79756 157150 79908
rect 157288 79840 157294 79892
rect 157346 79840 157352 79892
rect 157122 79716 157156 79756
rect 157150 79704 157156 79716
rect 157208 79704 157214 79756
rect 157306 79688 157334 79840
rect 157242 79636 157248 79688
rect 157300 79648 157334 79688
rect 157300 79636 157306 79648
rect 157398 79620 157426 79908
rect 157334 79568 157340 79620
rect 157392 79580 157426 79620
rect 157490 79620 157518 79908
rect 157582 79688 157610 79908
rect 157840 79880 157846 79892
rect 157766 79852 157846 79880
rect 157766 79744 157794 79852
rect 157840 79840 157846 79852
rect 157898 79840 157904 79892
rect 157720 79716 157794 79744
rect 157582 79648 157616 79688
rect 157610 79636 157616 79648
rect 157668 79636 157674 79688
rect 157490 79580 157524 79620
rect 157392 79568 157398 79580
rect 157518 79568 157524 79580
rect 157576 79568 157582 79620
rect 156656 79512 156920 79540
rect 156656 79500 156662 79512
rect 157058 79500 157064 79552
rect 157116 79540 157122 79552
rect 157720 79540 157748 79716
rect 157794 79568 157800 79620
rect 157852 79608 157858 79620
rect 157950 79608 157978 79920
rect 158300 79908 158306 79960
rect 158358 79908 158364 79960
rect 158392 79908 158398 79960
rect 158450 79908 158456 79960
rect 158576 79908 158582 79960
rect 158634 79908 158640 79960
rect 158668 79908 158674 79960
rect 158726 79908 158732 79960
rect 159128 79908 159134 79960
rect 159186 79908 159192 79960
rect 159220 79908 159226 79960
rect 159278 79908 159284 79960
rect 159496 79908 159502 79960
rect 159554 79908 159560 79960
rect 159680 79908 159686 79960
rect 159738 79908 159744 79960
rect 159772 79908 159778 79960
rect 159830 79908 159836 79960
rect 160048 79908 160054 79960
rect 160106 79908 160112 79960
rect 160140 79908 160146 79960
rect 160198 79908 160204 79960
rect 160232 79908 160238 79960
rect 160290 79908 160296 79960
rect 160416 79908 160422 79960
rect 160474 79908 160480 79960
rect 160600 79908 160606 79960
rect 160658 79908 160664 79960
rect 160784 79908 160790 79960
rect 160842 79908 160848 79960
rect 160876 79908 160882 79960
rect 160934 79908 160940 79960
rect 161244 79908 161250 79960
rect 161302 79908 161308 79960
rect 161428 79908 161434 79960
rect 161486 79908 161492 79960
rect 161704 79908 161710 79960
rect 161762 79908 161768 79960
rect 162072 79908 162078 79960
rect 162130 79908 162136 79960
rect 158024 79840 158030 79892
rect 158082 79840 158088 79892
rect 158208 79840 158214 79892
rect 158266 79840 158272 79892
rect 157852 79580 157978 79608
rect 157852 79568 157858 79580
rect 158042 79552 158070 79840
rect 158116 79772 158122 79824
rect 158174 79772 158180 79824
rect 158134 79688 158162 79772
rect 158226 79756 158254 79840
rect 158318 79824 158346 79908
rect 158410 79880 158438 79908
rect 158410 79852 158484 79880
rect 158456 79824 158484 79852
rect 158594 79824 158622 79908
rect 158318 79784 158352 79824
rect 158346 79772 158352 79784
rect 158404 79772 158410 79824
rect 158438 79772 158444 79824
rect 158496 79772 158502 79824
rect 158576 79772 158582 79824
rect 158634 79772 158640 79824
rect 158226 79716 158260 79756
rect 158254 79704 158260 79716
rect 158312 79704 158318 79756
rect 158686 79688 158714 79908
rect 158852 79840 158858 79892
rect 158910 79840 158916 79892
rect 158944 79840 158950 79892
rect 159002 79840 159008 79892
rect 158134 79648 158168 79688
rect 158162 79636 158168 79648
rect 158220 79636 158226 79688
rect 158622 79636 158628 79688
rect 158680 79648 158714 79688
rect 158680 79636 158686 79648
rect 157116 79512 157748 79540
rect 157116 79500 157122 79512
rect 157978 79500 157984 79552
rect 158036 79512 158070 79552
rect 158870 79552 158898 79840
rect 158962 79620 158990 79840
rect 159146 79688 159174 79908
rect 159238 79744 159266 79908
rect 159514 79744 159542 79908
rect 159238 79716 159312 79744
rect 159146 79648 159180 79688
rect 159174 79636 159180 79648
rect 159232 79636 159238 79688
rect 158962 79580 158996 79620
rect 158990 79568 158996 79580
rect 159048 79568 159054 79620
rect 159082 79568 159088 79620
rect 159140 79608 159146 79620
rect 159284 79608 159312 79716
rect 159140 79580 159312 79608
rect 159376 79716 159542 79744
rect 159140 79568 159146 79580
rect 158870 79512 158904 79552
rect 158036 79500 158042 79512
rect 158898 79500 158904 79512
rect 158956 79500 158962 79552
rect 159266 79500 159272 79552
rect 159324 79540 159330 79552
rect 159376 79540 159404 79716
rect 159542 79568 159548 79620
rect 159600 79608 159606 79620
rect 159698 79608 159726 79908
rect 159600 79580 159726 79608
rect 159790 79620 159818 79908
rect 160066 79812 160094 79908
rect 160020 79784 160094 79812
rect 159790 79580 159824 79620
rect 159600 79568 159606 79580
rect 159818 79568 159824 79580
rect 159876 79568 159882 79620
rect 159324 79512 159404 79540
rect 159324 79500 159330 79512
rect 153068 79444 153424 79472
rect 153068 79432 153074 79444
rect 154206 79432 154212 79484
rect 154264 79472 154270 79484
rect 158346 79472 158352 79484
rect 154264 79444 158352 79472
rect 154264 79432 154270 79444
rect 158346 79432 158352 79444
rect 158404 79432 158410 79484
rect 158622 79432 158628 79484
rect 158680 79472 158686 79484
rect 160020 79472 160048 79784
rect 160158 79744 160186 79908
rect 160112 79716 160186 79744
rect 160112 79540 160140 79716
rect 160250 79688 160278 79908
rect 160324 79840 160330 79892
rect 160382 79840 160388 79892
rect 160186 79636 160192 79688
rect 160244 79648 160278 79688
rect 160244 79636 160250 79648
rect 160342 79608 160370 79840
rect 160434 79824 160462 79908
rect 160434 79784 160468 79824
rect 160462 79772 160468 79784
rect 160520 79772 160526 79824
rect 160618 79756 160646 79908
rect 160554 79704 160560 79756
rect 160612 79716 160646 79756
rect 160612 79704 160618 79716
rect 160802 79688 160830 79908
rect 160738 79636 160744 79688
rect 160796 79648 160830 79688
rect 160796 79636 160802 79648
rect 160894 79620 160922 79908
rect 161060 79880 161066 79892
rect 160342 79580 160508 79608
rect 160480 79552 160508 79580
rect 160830 79568 160836 79620
rect 160888 79580 160922 79620
rect 160986 79852 161066 79880
rect 160888 79568 160894 79580
rect 160986 79552 161014 79852
rect 161060 79840 161066 79852
rect 161118 79840 161124 79892
rect 161152 79840 161158 79892
rect 161210 79840 161216 79892
rect 161170 79552 161198 79840
rect 161262 79756 161290 79908
rect 161262 79716 161296 79756
rect 161290 79704 161296 79716
rect 161348 79704 161354 79756
rect 160278 79540 160284 79552
rect 160112 79512 160284 79540
rect 160278 79500 160284 79512
rect 160336 79500 160342 79552
rect 160462 79500 160468 79552
rect 160520 79500 160526 79552
rect 160922 79500 160928 79552
rect 160980 79512 161014 79552
rect 160980 79500 160986 79512
rect 161106 79500 161112 79552
rect 161164 79512 161198 79552
rect 161446 79540 161474 79908
rect 161888 79840 161894 79892
rect 161946 79840 161952 79892
rect 162090 79880 162118 79908
rect 162090 79852 162210 79880
rect 161796 79812 161802 79824
rect 161768 79772 161802 79812
rect 161854 79772 161860 79824
rect 161906 79812 161934 79840
rect 161906 79784 162072 79812
rect 161658 79704 161664 79756
rect 161716 79744 161722 79756
rect 161768 79744 161796 79772
rect 161716 79716 161796 79744
rect 161716 79704 161722 79716
rect 162044 79552 162072 79784
rect 162182 79744 162210 79852
rect 162256 79772 162262 79824
rect 162314 79812 162320 79824
rect 162314 79772 162348 79812
rect 162182 79716 162256 79744
rect 162228 79620 162256 79716
rect 162210 79568 162216 79620
rect 162268 79568 162274 79620
rect 161566 79540 161572 79552
rect 161446 79512 161572 79540
rect 161164 79500 161170 79512
rect 161566 79500 161572 79512
rect 161624 79500 161630 79552
rect 162026 79500 162032 79552
rect 162084 79500 162090 79552
rect 158680 79444 160048 79472
rect 158680 79432 158686 79444
rect 161474 79432 161480 79484
rect 161532 79472 161538 79484
rect 162320 79472 162348 79772
rect 162412 79688 162440 79988
rect 164206 79988 168558 80016
rect 162532 79908 162538 79960
rect 162590 79908 162596 79960
rect 162808 79908 162814 79960
rect 162866 79908 162872 79960
rect 162900 79908 162906 79960
rect 162958 79908 162964 79960
rect 163820 79948 163826 79960
rect 163332 79920 163826 79948
rect 162394 79636 162400 79688
rect 162452 79636 162458 79688
rect 162550 79484 162578 79908
rect 162826 79824 162854 79908
rect 162808 79772 162814 79824
rect 162866 79772 162872 79824
rect 161532 79444 162348 79472
rect 161532 79432 161538 79444
rect 162486 79432 162492 79484
rect 162544 79444 162578 79484
rect 162544 79432 162550 79444
rect 162762 79432 162768 79484
rect 162820 79472 162826 79484
rect 162918 79472 162946 79908
rect 162992 79772 162998 79824
rect 163050 79772 163056 79824
rect 163010 79540 163038 79772
rect 163332 79608 163360 79920
rect 163820 79908 163826 79920
rect 163878 79908 163884 79960
rect 163912 79908 163918 79960
rect 163970 79908 163976 79960
rect 163452 79880 163458 79892
rect 163424 79840 163458 79880
rect 163510 79840 163516 79892
rect 163544 79840 163550 79892
rect 163602 79840 163608 79892
rect 163728 79840 163734 79892
rect 163786 79840 163792 79892
rect 163930 79880 163958 79908
rect 163884 79852 163958 79880
rect 163424 79676 163452 79840
rect 163562 79756 163590 79840
rect 163498 79704 163504 79756
rect 163556 79716 163590 79756
rect 163746 79744 163774 79840
rect 163700 79716 163774 79744
rect 163556 79704 163562 79716
rect 163700 79688 163728 79716
rect 163590 79676 163596 79688
rect 163424 79648 163596 79676
rect 163590 79636 163596 79648
rect 163648 79636 163654 79688
rect 163682 79636 163688 79688
rect 163740 79636 163746 79688
rect 163884 79620 163912 79852
rect 164004 79812 164010 79824
rect 163976 79772 164010 79812
rect 164062 79772 164068 79824
rect 163976 79688 164004 79772
rect 164206 79744 164234 79988
rect 164464 79908 164470 79960
rect 164522 79948 164528 79960
rect 164522 79920 164694 79948
rect 164522 79908 164528 79920
rect 164280 79840 164286 79892
rect 164338 79840 164344 79892
rect 164556 79840 164562 79892
rect 164614 79840 164620 79892
rect 164114 79716 164234 79744
rect 164298 79756 164326 79840
rect 164298 79716 164332 79756
rect 163958 79636 163964 79688
rect 164016 79636 164022 79688
rect 164114 79676 164142 79716
rect 164326 79704 164332 79716
rect 164384 79704 164390 79756
rect 164574 79676 164602 79840
rect 164068 79648 164142 79676
rect 164344 79648 164602 79676
rect 164068 79620 164096 79648
rect 163774 79608 163780 79620
rect 163332 79580 163780 79608
rect 163774 79568 163780 79580
rect 163832 79568 163838 79620
rect 163866 79568 163872 79620
rect 163924 79568 163930 79620
rect 164050 79568 164056 79620
rect 164108 79568 164114 79620
rect 164234 79568 164240 79620
rect 164292 79608 164298 79620
rect 164344 79608 164372 79648
rect 164292 79580 164372 79608
rect 164292 79568 164298 79580
rect 164666 79552 164694 79920
rect 165752 79908 165758 79960
rect 165810 79948 165816 79960
rect 165936 79948 165942 79960
rect 165810 79908 165844 79948
rect 164924 79840 164930 79892
rect 164982 79840 164988 79892
rect 165016 79840 165022 79892
rect 165074 79840 165080 79892
rect 165108 79840 165114 79892
rect 165166 79880 165172 79892
rect 165166 79840 165200 79880
rect 165292 79840 165298 79892
rect 165350 79840 165356 79892
rect 165660 79840 165666 79892
rect 165718 79840 165724 79892
rect 164942 79756 164970 79840
rect 165034 79812 165062 79840
rect 165034 79784 165108 79812
rect 164942 79716 164976 79756
rect 164970 79704 164976 79716
rect 165028 79704 165034 79756
rect 165080 79688 165108 79784
rect 165172 79756 165200 79840
rect 165310 79756 165338 79840
rect 165568 79772 165574 79824
rect 165626 79772 165632 79824
rect 165154 79704 165160 79756
rect 165212 79704 165218 79756
rect 165246 79704 165252 79756
rect 165304 79716 165338 79756
rect 165304 79704 165310 79716
rect 165586 79688 165614 79772
rect 165678 79756 165706 79840
rect 165678 79716 165712 79756
rect 165706 79704 165712 79716
rect 165764 79704 165770 79756
rect 165816 79688 165844 79908
rect 165908 79908 165942 79948
rect 165994 79908 166000 79960
rect 166028 79908 166034 79960
rect 166086 79908 166092 79960
rect 166120 79908 166126 79960
rect 166178 79908 166184 79960
rect 166856 79948 166862 79960
rect 166506 79920 166862 79948
rect 165062 79636 165068 79688
rect 165120 79636 165126 79688
rect 165522 79636 165528 79688
rect 165580 79648 165614 79688
rect 165580 79636 165586 79648
rect 165798 79636 165804 79688
rect 165856 79636 165862 79688
rect 165908 79676 165936 79908
rect 166046 79880 166074 79908
rect 166000 79852 166074 79880
rect 166000 79824 166028 79852
rect 166138 79824 166166 79908
rect 166396 79840 166402 79892
rect 166454 79840 166460 79892
rect 165982 79772 165988 79824
rect 166040 79772 166046 79824
rect 166074 79772 166080 79824
rect 166132 79784 166166 79824
rect 166132 79772 166138 79784
rect 166212 79772 166218 79824
rect 166270 79812 166276 79824
rect 166270 79772 166304 79812
rect 166166 79676 166172 79688
rect 165908 79648 166172 79676
rect 166166 79636 166172 79648
rect 166224 79636 166230 79688
rect 165982 79568 165988 79620
rect 166040 79568 166046 79620
rect 164418 79540 164424 79552
rect 163010 79512 164424 79540
rect 164418 79500 164424 79512
rect 164476 79500 164482 79552
rect 164666 79512 164700 79552
rect 164694 79500 164700 79512
rect 164752 79500 164758 79552
rect 162820 79444 162946 79472
rect 162820 79432 162826 79444
rect 163038 79432 163044 79484
rect 163096 79472 163102 79484
rect 163498 79472 163504 79484
rect 163096 79444 163504 79472
rect 163096 79432 163102 79444
rect 163498 79432 163504 79444
rect 163556 79432 163562 79484
rect 152642 79404 152648 79416
rect 150360 79376 152648 79404
rect 152642 79364 152648 79376
rect 152700 79364 152706 79416
rect 158070 79404 158076 79416
rect 153764 79376 158076 79404
rect 3970 79296 3976 79348
rect 4028 79336 4034 79348
rect 4028 79308 140268 79336
rect 4028 79296 4034 79308
rect 130194 79228 130200 79280
rect 130252 79268 130258 79280
rect 132678 79268 132684 79280
rect 130252 79240 132684 79268
rect 130252 79228 130258 79240
rect 132678 79228 132684 79240
rect 132736 79228 132742 79280
rect 134518 79228 134524 79280
rect 134576 79268 134582 79280
rect 140130 79268 140136 79280
rect 134576 79240 140136 79268
rect 134576 79228 134582 79240
rect 140130 79228 140136 79240
rect 140188 79228 140194 79280
rect 129366 79160 129372 79212
rect 129424 79200 129430 79212
rect 140038 79200 140044 79212
rect 129424 79172 140044 79200
rect 129424 79160 129430 79172
rect 140038 79160 140044 79172
rect 140096 79160 140102 79212
rect 137278 79092 137284 79144
rect 137336 79132 137342 79144
rect 140130 79132 140136 79144
rect 137336 79104 140136 79132
rect 137336 79092 137342 79104
rect 140130 79092 140136 79104
rect 140188 79092 140194 79144
rect 140240 79132 140268 79308
rect 140958 79296 140964 79348
rect 141016 79336 141022 79348
rect 141970 79336 141976 79348
rect 141016 79308 141976 79336
rect 141016 79296 141022 79308
rect 141970 79296 141976 79308
rect 142028 79296 142034 79348
rect 149238 79296 149244 79348
rect 149296 79336 149302 79348
rect 153764 79336 153792 79376
rect 158070 79364 158076 79376
rect 158128 79364 158134 79416
rect 158530 79364 158536 79416
rect 158588 79404 158594 79416
rect 165614 79404 165620 79416
rect 158588 79376 165620 79404
rect 158588 79364 158594 79376
rect 165614 79364 165620 79376
rect 165672 79364 165678 79416
rect 165890 79364 165896 79416
rect 165948 79404 165954 79416
rect 166000 79404 166028 79568
rect 165948 79376 166028 79404
rect 166276 79404 166304 79772
rect 166414 79676 166442 79840
rect 166368 79648 166442 79676
rect 166368 79484 166396 79648
rect 166350 79432 166356 79484
rect 166408 79432 166414 79484
rect 166506 79472 166534 79920
rect 166856 79908 166862 79920
rect 166914 79908 166920 79960
rect 167132 79948 167138 79960
rect 167058 79920 167138 79948
rect 166764 79840 166770 79892
rect 166822 79840 166828 79892
rect 166948 79840 166954 79892
rect 167006 79840 167012 79892
rect 166782 79620 166810 79840
rect 166782 79580 166816 79620
rect 166810 79568 166816 79580
rect 166868 79568 166874 79620
rect 166626 79500 166632 79552
rect 166684 79540 166690 79552
rect 166966 79540 166994 79840
rect 167058 79756 167086 79920
rect 167132 79908 167138 79920
rect 167190 79908 167196 79960
rect 167592 79908 167598 79960
rect 167650 79908 167656 79960
rect 167776 79948 167782 79960
rect 167702 79920 167782 79948
rect 167224 79880 167230 79892
rect 167196 79840 167230 79880
rect 167282 79840 167288 79892
rect 167408 79840 167414 79892
rect 167466 79840 167472 79892
rect 167610 79880 167638 79908
rect 167564 79852 167638 79880
rect 167702 79880 167730 79920
rect 167776 79908 167782 79920
rect 167834 79908 167840 79960
rect 167868 79908 167874 79960
rect 167926 79908 167932 79960
rect 167960 79908 167966 79960
rect 168018 79908 168024 79960
rect 168052 79908 168058 79960
rect 168110 79908 168116 79960
rect 167886 79880 167914 79908
rect 167702 79852 167776 79880
rect 167196 79756 167224 79840
rect 167426 79756 167454 79840
rect 167058 79716 167092 79756
rect 167086 79704 167092 79716
rect 167144 79704 167150 79756
rect 167178 79704 167184 79756
rect 167236 79704 167242 79756
rect 167426 79716 167460 79756
rect 167454 79704 167460 79716
rect 167512 79704 167518 79756
rect 167564 79688 167592 79852
rect 167546 79636 167552 79688
rect 167604 79636 167610 79688
rect 167748 79620 167776 79852
rect 167840 79852 167914 79880
rect 167840 79620 167868 79852
rect 167978 79756 168006 79908
rect 167914 79704 167920 79756
rect 167972 79716 168006 79756
rect 167972 79704 167978 79716
rect 167730 79568 167736 79620
rect 167788 79568 167794 79620
rect 167822 79568 167828 79620
rect 167880 79568 167886 79620
rect 168070 79608 168098 79908
rect 168530 79676 168558 79988
rect 169450 79988 169662 80016
rect 170462 79988 172514 80016
rect 172946 79988 173434 80016
rect 169450 79960 169478 79988
rect 168788 79908 168794 79960
rect 168846 79908 168852 79960
rect 169432 79908 169438 79960
rect 169490 79908 169496 79960
rect 168604 79840 168610 79892
rect 168662 79840 168668 79892
rect 168622 79756 168650 79840
rect 168622 79716 168656 79756
rect 168650 79704 168656 79716
rect 168708 79704 168714 79756
rect 168530 79648 168650 79676
rect 168282 79608 168288 79620
rect 168070 79580 168288 79608
rect 168282 79568 168288 79580
rect 168340 79568 168346 79620
rect 166684 79512 166994 79540
rect 166684 79500 166690 79512
rect 166902 79472 166908 79484
rect 166506 79444 166908 79472
rect 166902 79432 166908 79444
rect 166960 79432 166966 79484
rect 168098 79432 168104 79484
rect 168156 79472 168162 79484
rect 168622 79472 168650 79648
rect 168806 79608 168834 79908
rect 168880 79840 168886 79892
rect 168938 79840 168944 79892
rect 169340 79880 169346 79892
rect 169312 79840 169346 79880
rect 169398 79840 169404 79892
rect 169524 79840 169530 79892
rect 169582 79840 169588 79892
rect 168898 79744 168926 79840
rect 168898 79716 169156 79744
rect 169018 79608 169024 79620
rect 168806 79580 169024 79608
rect 169018 79568 169024 79580
rect 169076 79568 169082 79620
rect 168834 79500 168840 79552
rect 168892 79540 168898 79552
rect 169128 79540 169156 79716
rect 169312 79620 169340 79840
rect 169386 79704 169392 79756
rect 169444 79744 169450 79756
rect 169542 79744 169570 79840
rect 169444 79716 169570 79744
rect 169444 79704 169450 79716
rect 169478 79636 169484 79688
rect 169536 79676 169542 79688
rect 169634 79676 169662 79988
rect 172946 79960 172974 79988
rect 169800 79908 169806 79960
rect 169858 79908 169864 79960
rect 169892 79908 169898 79960
rect 169950 79908 169956 79960
rect 169984 79908 169990 79960
rect 170042 79908 170048 79960
rect 170168 79908 170174 79960
rect 170226 79908 170232 79960
rect 170812 79908 170818 79960
rect 170870 79908 170876 79960
rect 171548 79908 171554 79960
rect 171606 79908 171612 79960
rect 171640 79908 171646 79960
rect 171698 79948 171704 79960
rect 171824 79948 171830 79960
rect 171698 79908 171732 79948
rect 169818 79756 169846 79908
rect 169754 79704 169760 79756
rect 169812 79716 169846 79756
rect 169812 79704 169818 79716
rect 169536 79648 169662 79676
rect 169536 79636 169542 79648
rect 169294 79568 169300 79620
rect 169352 79568 169358 79620
rect 168892 79512 169156 79540
rect 168892 79500 168898 79512
rect 169910 79472 169938 79908
rect 170002 79688 170030 79908
rect 170186 79756 170214 79908
rect 170444 79840 170450 79892
rect 170502 79840 170508 79892
rect 170536 79840 170542 79892
rect 170594 79880 170600 79892
rect 170594 79840 170628 79880
rect 170122 79704 170128 79756
rect 170180 79716 170214 79756
rect 170462 79756 170490 79840
rect 170462 79716 170496 79756
rect 170180 79704 170186 79716
rect 170490 79704 170496 79716
rect 170548 79704 170554 79756
rect 170002 79648 170036 79688
rect 170030 79636 170036 79648
rect 170088 79636 170094 79688
rect 170030 79500 170036 79552
rect 170088 79540 170094 79552
rect 170600 79540 170628 79840
rect 170674 79636 170680 79688
rect 170732 79676 170738 79688
rect 170830 79676 170858 79908
rect 171364 79880 171370 79892
rect 171336 79840 171370 79880
rect 171422 79840 171428 79892
rect 171336 79756 171364 79840
rect 171318 79704 171324 79756
rect 171376 79704 171382 79756
rect 170732 79648 170858 79676
rect 171566 79688 171594 79908
rect 171566 79648 171600 79688
rect 170732 79636 170738 79648
rect 171594 79636 171600 79648
rect 171652 79636 171658 79688
rect 170088 79512 170628 79540
rect 170088 79500 170094 79512
rect 171226 79500 171232 79552
rect 171284 79540 171290 79552
rect 171704 79540 171732 79908
rect 171796 79908 171830 79948
rect 171882 79908 171888 79960
rect 171916 79908 171922 79960
rect 171974 79908 171980 79960
rect 172008 79908 172014 79960
rect 172066 79908 172072 79960
rect 172468 79908 172474 79960
rect 172526 79908 172532 79960
rect 172560 79908 172566 79960
rect 172618 79908 172624 79960
rect 172744 79908 172750 79960
rect 172802 79908 172808 79960
rect 172928 79908 172934 79960
rect 172986 79908 172992 79960
rect 173112 79908 173118 79960
rect 173170 79908 173176 79960
rect 171796 79756 171824 79908
rect 171778 79704 171784 79756
rect 171836 79704 171842 79756
rect 171284 79512 171732 79540
rect 171284 79500 171290 79512
rect 170306 79472 170312 79484
rect 168156 79444 168374 79472
rect 168622 79444 169708 79472
rect 169910 79444 170312 79472
rect 168156 79432 168162 79444
rect 166626 79404 166632 79416
rect 166276 79376 166632 79404
rect 165948 79364 165954 79376
rect 166626 79364 166632 79376
rect 166684 79364 166690 79416
rect 166994 79364 167000 79416
rect 167052 79404 167058 79416
rect 167270 79404 167276 79416
rect 167052 79376 167276 79404
rect 167052 79364 167058 79376
rect 167270 79364 167276 79376
rect 167328 79364 167334 79416
rect 168346 79404 168374 79444
rect 168558 79404 168564 79416
rect 168346 79376 168564 79404
rect 168558 79364 168564 79376
rect 168616 79364 168622 79416
rect 169570 79336 169576 79348
rect 149296 79308 153792 79336
rect 153856 79308 169576 79336
rect 149296 79296 149302 79308
rect 153856 79268 153884 79308
rect 169570 79296 169576 79308
rect 169628 79296 169634 79348
rect 169680 79336 169708 79444
rect 170306 79432 170312 79444
rect 170364 79432 170370 79484
rect 171410 79432 171416 79484
rect 171468 79472 171474 79484
rect 171934 79472 171962 79908
rect 172026 79824 172054 79908
rect 172192 79840 172198 79892
rect 172250 79840 172256 79892
rect 172008 79772 172014 79824
rect 172066 79772 172072 79824
rect 172100 79772 172106 79824
rect 172158 79772 172164 79824
rect 172118 79620 172146 79772
rect 172054 79568 172060 79620
rect 172112 79580 172146 79620
rect 172112 79568 172118 79580
rect 172210 79552 172238 79840
rect 172284 79772 172290 79824
rect 172342 79772 172348 79824
rect 172486 79812 172514 79908
rect 172394 79784 172514 79812
rect 172146 79500 172152 79552
rect 172204 79512 172238 79552
rect 172204 79500 172210 79512
rect 172302 79484 172330 79772
rect 171468 79444 171962 79472
rect 171468 79432 171474 79444
rect 172238 79432 172244 79484
rect 172296 79444 172330 79484
rect 172296 79432 172302 79444
rect 172394 79416 172422 79784
rect 172578 79608 172606 79908
rect 170122 79364 170128 79416
rect 170180 79404 170186 79416
rect 170490 79404 170496 79416
rect 170180 79376 170496 79404
rect 170180 79364 170186 79376
rect 170490 79364 170496 79376
rect 170548 79364 170554 79416
rect 172330 79364 172336 79416
rect 172388 79376 172422 79416
rect 172532 79580 172606 79608
rect 172532 79404 172560 79580
rect 172606 79500 172612 79552
rect 172664 79540 172670 79552
rect 172762 79540 172790 79908
rect 173130 79880 173158 79908
rect 172946 79852 173158 79880
rect 172946 79744 172974 79852
rect 173296 79840 173302 79892
rect 173354 79840 173360 79892
rect 173020 79772 173026 79824
rect 173078 79772 173084 79824
rect 172900 79716 172974 79744
rect 172900 79676 172928 79716
rect 173038 79688 173066 79772
rect 172664 79512 172790 79540
rect 172854 79648 172928 79676
rect 172664 79500 172670 79512
rect 172698 79432 172704 79484
rect 172756 79472 172762 79484
rect 172854 79472 172882 79648
rect 172974 79636 172980 79688
rect 173032 79648 173066 79688
rect 173032 79636 173038 79648
rect 173314 79552 173342 79840
rect 173406 79620 173434 79988
rect 174050 79988 174446 80016
rect 174878 79988 175090 80016
rect 176902 79988 178126 80016
rect 173480 79908 173486 79960
rect 173538 79908 173544 79960
rect 173572 79908 173578 79960
rect 173630 79908 173636 79960
rect 173664 79908 173670 79960
rect 173722 79908 173728 79960
rect 173848 79908 173854 79960
rect 173906 79908 173912 79960
rect 173498 79688 173526 79908
rect 173590 79824 173618 79908
rect 173572 79772 173578 79824
rect 173630 79772 173636 79824
rect 173682 79688 173710 79908
rect 173498 79648 173532 79688
rect 173526 79636 173532 79648
rect 173584 79636 173590 79688
rect 173618 79636 173624 79688
rect 173676 79648 173710 79688
rect 173676 79636 173682 79648
rect 173406 79580 173440 79620
rect 173434 79568 173440 79580
rect 173492 79568 173498 79620
rect 173250 79500 173256 79552
rect 173308 79512 173342 79552
rect 173308 79500 173314 79512
rect 173710 79500 173716 79552
rect 173768 79540 173774 79552
rect 173866 79540 173894 79908
rect 173768 79512 173894 79540
rect 174050 79552 174078 79988
rect 174418 79960 174446 79988
rect 176902 79960 176930 79988
rect 174216 79908 174222 79960
rect 174274 79908 174280 79960
rect 174308 79908 174314 79960
rect 174366 79908 174372 79960
rect 174400 79908 174406 79960
rect 174458 79908 174464 79960
rect 174492 79908 174498 79960
rect 174550 79908 174556 79960
rect 174584 79908 174590 79960
rect 174642 79908 174648 79960
rect 174768 79908 174774 79960
rect 174826 79908 174832 79960
rect 174860 79908 174866 79960
rect 174918 79908 174924 79960
rect 175044 79908 175050 79960
rect 175102 79908 175108 79960
rect 175320 79908 175326 79960
rect 175378 79908 175384 79960
rect 175964 79908 175970 79960
rect 176022 79908 176028 79960
rect 176148 79908 176154 79960
rect 176206 79908 176212 79960
rect 176332 79908 176338 79960
rect 176390 79948 176396 79960
rect 176390 79908 176424 79948
rect 176516 79908 176522 79960
rect 176574 79908 176580 79960
rect 176608 79908 176614 79960
rect 176666 79908 176672 79960
rect 176700 79908 176706 79960
rect 176758 79908 176764 79960
rect 176792 79908 176798 79960
rect 176850 79908 176856 79960
rect 176884 79908 176890 79960
rect 176942 79908 176948 79960
rect 176976 79908 176982 79960
rect 177034 79908 177040 79960
rect 177068 79908 177074 79960
rect 177126 79908 177132 79960
rect 177252 79948 177258 79960
rect 177178 79920 177258 79948
rect 174050 79512 174084 79552
rect 173768 79500 173774 79512
rect 174078 79500 174084 79512
rect 174136 79500 174142 79552
rect 174234 79540 174262 79908
rect 174326 79608 174354 79908
rect 174510 79756 174538 79908
rect 174446 79704 174452 79756
rect 174504 79716 174538 79756
rect 174504 79704 174510 79716
rect 174602 79676 174630 79908
rect 174786 79824 174814 79908
rect 174768 79772 174774 79824
rect 174826 79772 174832 79824
rect 174878 79676 174906 79908
rect 175062 79756 175090 79908
rect 175136 79840 175142 79892
rect 175194 79880 175200 79892
rect 175194 79840 175228 79880
rect 175200 79756 175228 79840
rect 175062 79716 175096 79756
rect 175090 79704 175096 79716
rect 175148 79704 175154 79756
rect 175182 79704 175188 79756
rect 175240 79704 175246 79756
rect 175338 79688 175366 79908
rect 175982 79756 176010 79908
rect 176056 79840 176062 79892
rect 176114 79840 176120 79892
rect 176166 79880 176194 79908
rect 176166 79852 176332 79880
rect 176074 79812 176102 79840
rect 176074 79784 176148 79812
rect 176120 79756 176148 79784
rect 175982 79716 176016 79756
rect 176010 79704 176016 79716
rect 176068 79704 176074 79756
rect 176102 79704 176108 79756
rect 176160 79704 176166 79756
rect 174602 79648 174676 79676
rect 174878 79648 175044 79676
rect 175338 79648 175372 79688
rect 174538 79608 174544 79620
rect 174326 79580 174544 79608
rect 174538 79568 174544 79580
rect 174596 79568 174602 79620
rect 174446 79540 174452 79552
rect 174234 79512 174452 79540
rect 174446 79500 174452 79512
rect 174504 79500 174510 79552
rect 172756 79444 172882 79472
rect 172756 79432 172762 79444
rect 174538 79432 174544 79484
rect 174596 79472 174602 79484
rect 174648 79472 174676 79648
rect 174722 79500 174728 79552
rect 174780 79540 174786 79552
rect 175016 79540 175044 79648
rect 175366 79636 175372 79648
rect 175424 79636 175430 79688
rect 174780 79512 175044 79540
rect 174780 79500 174786 79512
rect 174596 79444 174676 79472
rect 174596 79432 174602 79444
rect 172790 79404 172796 79416
rect 172532 79376 172796 79404
rect 172388 79364 172394 79376
rect 172790 79364 172796 79376
rect 172848 79364 172854 79416
rect 173158 79364 173164 79416
rect 173216 79404 173222 79416
rect 175458 79404 175464 79416
rect 173216 79376 175464 79404
rect 173216 79364 173222 79376
rect 175458 79364 175464 79376
rect 175516 79364 175522 79416
rect 176304 79404 176332 79852
rect 176396 79688 176424 79908
rect 176534 79880 176562 79908
rect 176488 79852 176562 79880
rect 176488 79756 176516 79852
rect 176626 79756 176654 79908
rect 176470 79704 176476 79756
rect 176528 79704 176534 79756
rect 176562 79704 176568 79756
rect 176620 79716 176654 79756
rect 176620 79704 176626 79716
rect 176378 79636 176384 79688
rect 176436 79636 176442 79688
rect 176718 79676 176746 79908
rect 176810 79756 176838 79908
rect 176994 79756 177022 79908
rect 176810 79716 176844 79756
rect 176838 79704 176844 79716
rect 176896 79704 176902 79756
rect 176930 79704 176936 79756
rect 176988 79716 177022 79756
rect 176988 79704 176994 79716
rect 176718 79648 176792 79676
rect 176764 79472 176792 79648
rect 176838 79500 176844 79552
rect 176896 79540 176902 79552
rect 177086 79540 177114 79908
rect 177178 79756 177206 79920
rect 177252 79908 177258 79920
rect 177310 79908 177316 79960
rect 177344 79908 177350 79960
rect 177402 79908 177408 79960
rect 178098 79948 178126 79988
rect 178466 79960 178494 80056
rect 188890 80044 188896 80096
rect 188948 80084 188954 80096
rect 580442 80084 580448 80096
rect 188948 80056 580448 80084
rect 188948 80044 188954 80056
rect 580442 80044 580448 80056
rect 580500 80044 580506 80096
rect 178926 79988 179552 80016
rect 178926 79960 178954 79988
rect 178098 79920 178172 79948
rect 177362 79880 177390 79908
rect 177316 79852 177390 79880
rect 177316 79824 177344 79852
rect 177436 79840 177442 79892
rect 177494 79840 177500 79892
rect 177712 79840 177718 79892
rect 177770 79880 177776 79892
rect 177770 79852 178080 79880
rect 177770 79840 177776 79852
rect 177298 79772 177304 79824
rect 177356 79772 177362 79824
rect 177178 79716 177212 79756
rect 177206 79704 177212 79716
rect 177264 79704 177270 79756
rect 176896 79512 177114 79540
rect 177454 79540 177482 79840
rect 177804 79772 177810 79824
rect 177862 79812 177868 79824
rect 177862 79772 177896 79812
rect 177868 79744 177896 79772
rect 178052 79744 178080 79852
rect 178144 79812 178172 79920
rect 178448 79908 178454 79960
rect 178506 79908 178512 79960
rect 178908 79908 178914 79960
rect 178966 79908 178972 79960
rect 179524 79948 179552 79988
rect 179966 79976 179972 80028
rect 180024 80016 180030 80028
rect 180024 79988 186314 80016
rect 180024 79976 180030 79988
rect 179690 79948 179696 79960
rect 179524 79920 179696 79948
rect 179690 79908 179696 79920
rect 179748 79908 179754 79960
rect 179276 79840 179282 79892
rect 179334 79880 179340 79892
rect 179782 79880 179788 79892
rect 179334 79852 179788 79880
rect 179334 79840 179340 79852
rect 179782 79840 179788 79852
rect 179840 79840 179846 79892
rect 180242 79812 180248 79824
rect 178144 79784 180248 79812
rect 180242 79772 180248 79784
rect 180300 79772 180306 79824
rect 186286 79812 186314 79988
rect 194226 79812 194232 79824
rect 186286 79784 194232 79812
rect 194226 79772 194232 79784
rect 194284 79772 194290 79824
rect 180518 79744 180524 79756
rect 177868 79716 177988 79744
rect 178052 79716 180524 79744
rect 177960 79608 177988 79716
rect 180518 79704 180524 79716
rect 180576 79704 180582 79756
rect 181714 79608 181720 79620
rect 177960 79580 181720 79608
rect 181714 79568 181720 79580
rect 181772 79568 181778 79620
rect 415394 79540 415400 79552
rect 177454 79512 177620 79540
rect 176896 79500 176902 79512
rect 177390 79472 177396 79484
rect 176764 79444 177396 79472
rect 177390 79432 177396 79444
rect 177448 79432 177454 79484
rect 177592 79472 177620 79512
rect 186286 79512 415400 79540
rect 178034 79472 178040 79484
rect 177592 79444 178040 79472
rect 178034 79432 178040 79444
rect 178092 79432 178098 79484
rect 178126 79432 178132 79484
rect 178184 79472 178190 79484
rect 186286 79472 186314 79512
rect 415394 79500 415400 79512
rect 415452 79500 415458 79552
rect 178184 79444 186314 79472
rect 178184 79432 178190 79444
rect 189718 79404 189724 79416
rect 176304 79376 189724 79404
rect 189718 79364 189724 79376
rect 189776 79364 189782 79416
rect 173066 79336 173072 79348
rect 169680 79308 173072 79336
rect 173066 79296 173072 79308
rect 173124 79296 173130 79348
rect 176746 79336 176752 79348
rect 173176 79308 176752 79336
rect 173176 79268 173204 79308
rect 176746 79296 176752 79308
rect 176804 79296 176810 79348
rect 177114 79296 177120 79348
rect 177172 79336 177178 79348
rect 179966 79336 179972 79348
rect 177172 79308 179972 79336
rect 177172 79296 177178 79308
rect 179966 79296 179972 79308
rect 180024 79296 180030 79348
rect 527174 79336 527180 79348
rect 180444 79308 527180 79336
rect 140746 79240 153884 79268
rect 154546 79240 173204 79268
rect 140746 79132 140774 79240
rect 140958 79160 140964 79212
rect 141016 79200 141022 79212
rect 141878 79200 141884 79212
rect 141016 79172 141884 79200
rect 141016 79160 141022 79172
rect 141878 79160 141884 79172
rect 141936 79160 141942 79212
rect 144454 79160 144460 79212
rect 144512 79200 144518 79212
rect 154546 79200 154574 79240
rect 173342 79228 173348 79280
rect 173400 79268 173406 79280
rect 174998 79268 175004 79280
rect 173400 79240 175004 79268
rect 173400 79228 173406 79240
rect 174998 79228 175004 79240
rect 175056 79228 175062 79280
rect 176378 79228 176384 79280
rect 176436 79268 176442 79280
rect 179874 79268 179880 79280
rect 176436 79240 179880 79268
rect 176436 79228 176442 79240
rect 179874 79228 179880 79240
rect 179932 79228 179938 79280
rect 144512 79172 154574 79200
rect 144512 79160 144518 79172
rect 157426 79160 157432 79212
rect 157484 79200 157490 79212
rect 159358 79200 159364 79212
rect 157484 79172 159364 79200
rect 157484 79160 157490 79172
rect 159358 79160 159364 79172
rect 159416 79160 159422 79212
rect 160094 79160 160100 79212
rect 160152 79200 160158 79212
rect 160152 79172 165752 79200
rect 160152 79160 160158 79172
rect 140240 79104 140774 79132
rect 158070 79092 158076 79144
rect 158128 79132 158134 79144
rect 164050 79132 164056 79144
rect 158128 79104 164056 79132
rect 158128 79092 158134 79104
rect 164050 79092 164056 79104
rect 164108 79092 164114 79144
rect 112438 79024 112444 79076
rect 112496 79064 112502 79076
rect 112496 79036 164234 79064
rect 112496 79024 112502 79036
rect 130010 78956 130016 79008
rect 130068 78996 130074 79008
rect 130838 78996 130844 79008
rect 130068 78968 130844 78996
rect 130068 78956 130074 78968
rect 130838 78956 130844 78968
rect 130896 78956 130902 79008
rect 137986 78968 157334 78996
rect 84838 78888 84844 78940
rect 84896 78928 84902 78940
rect 137986 78928 138014 78968
rect 84896 78900 138014 78928
rect 84896 78888 84902 78900
rect 140038 78888 140044 78940
rect 140096 78928 140102 78940
rect 144454 78928 144460 78940
rect 140096 78900 144460 78928
rect 140096 78888 140102 78900
rect 144454 78888 144460 78900
rect 144512 78888 144518 78940
rect 144914 78888 144920 78940
rect 144972 78928 144978 78940
rect 144972 78900 146800 78928
rect 144972 78888 144978 78900
rect 129366 78820 129372 78872
rect 129424 78860 129430 78872
rect 134150 78860 134156 78872
rect 129424 78832 134156 78860
rect 129424 78820 129430 78832
rect 134150 78820 134156 78832
rect 134208 78820 134214 78872
rect 135346 78820 135352 78872
rect 135404 78860 135410 78872
rect 146772 78860 146800 78900
rect 155310 78888 155316 78940
rect 155368 78888 155374 78940
rect 157306 78928 157334 78968
rect 158346 78956 158352 79008
rect 158404 78996 158410 79008
rect 160094 78996 160100 79008
rect 158404 78968 160100 78996
rect 158404 78956 158410 78968
rect 160094 78956 160100 78968
rect 160152 78956 160158 79008
rect 162578 78956 162584 79008
rect 162636 78996 162642 79008
rect 162854 78996 162860 79008
rect 162636 78968 162860 78996
rect 162636 78956 162642 78968
rect 162854 78956 162860 78968
rect 162912 78956 162918 79008
rect 163222 78956 163228 79008
rect 163280 78996 163286 79008
rect 163590 78996 163596 79008
rect 163280 78968 163596 78996
rect 163280 78956 163286 78968
rect 163590 78956 163596 78968
rect 163648 78956 163654 79008
rect 164206 78996 164234 79036
rect 164510 79024 164516 79076
rect 164568 79064 164574 79076
rect 164878 79064 164884 79076
rect 164568 79036 164884 79064
rect 164568 79024 164574 79036
rect 164878 79024 164884 79036
rect 164936 79024 164942 79076
rect 165724 79064 165752 79172
rect 165798 79160 165804 79212
rect 165856 79200 165862 79212
rect 176286 79200 176292 79212
rect 165856 79172 176292 79200
rect 165856 79160 165862 79172
rect 176286 79160 176292 79172
rect 176344 79160 176350 79212
rect 177298 79160 177304 79212
rect 177356 79200 177362 79212
rect 180444 79200 180472 79308
rect 527174 79296 527180 79308
rect 527232 79296 527238 79348
rect 180518 79228 180524 79280
rect 180576 79268 180582 79280
rect 192478 79268 192484 79280
rect 180576 79240 192484 79268
rect 180576 79228 180582 79240
rect 192478 79228 192484 79240
rect 192536 79228 192542 79280
rect 177356 79172 180472 79200
rect 177356 79160 177362 79172
rect 181714 79160 181720 79212
rect 181772 79200 181778 79212
rect 193858 79200 193864 79212
rect 181772 79172 193864 79200
rect 181772 79160 181778 79172
rect 193858 79160 193864 79172
rect 193916 79160 193922 79212
rect 166534 79092 166540 79144
rect 166592 79132 166598 79144
rect 171778 79132 171784 79144
rect 166592 79104 171784 79132
rect 166592 79092 166598 79104
rect 171778 79092 171784 79104
rect 171836 79092 171842 79144
rect 172422 79092 172428 79144
rect 172480 79132 172486 79144
rect 175274 79132 175280 79144
rect 172480 79104 175280 79132
rect 172480 79092 172486 79104
rect 175274 79092 175280 79104
rect 175332 79092 175338 79144
rect 178862 79132 178868 79144
rect 175384 79104 178868 79132
rect 168558 79064 168564 79076
rect 165724 79036 168564 79064
rect 168558 79024 168564 79036
rect 168616 79024 168622 79076
rect 169570 79024 169576 79076
rect 169628 79064 169634 79076
rect 175384 79064 175412 79104
rect 178862 79092 178868 79104
rect 178920 79092 178926 79144
rect 192662 79132 192668 79144
rect 186286 79104 192668 79132
rect 169628 79036 175412 79064
rect 169628 79024 169634 79036
rect 176654 79024 176660 79076
rect 176712 79064 176718 79076
rect 178126 79064 178132 79076
rect 176712 79036 178132 79064
rect 176712 79024 176718 79036
rect 178126 79024 178132 79036
rect 178184 79024 178190 79076
rect 179874 79024 179880 79076
rect 179932 79064 179938 79076
rect 186286 79064 186314 79104
rect 192662 79092 192668 79104
rect 192720 79092 192726 79144
rect 179932 79036 186314 79064
rect 179932 79024 179938 79036
rect 164206 78968 174492 78996
rect 170122 78928 170128 78940
rect 157306 78900 170128 78928
rect 170122 78888 170128 78900
rect 170180 78888 170186 78940
rect 170232 78900 171778 78928
rect 154206 78860 154212 78872
rect 135404 78832 140774 78860
rect 146772 78832 154212 78860
rect 135404 78820 135410 78832
rect 133874 78792 133880 78804
rect 125566 78764 133880 78792
rect 122098 78616 122104 78668
rect 122156 78656 122162 78668
rect 125566 78656 125594 78764
rect 133874 78752 133880 78764
rect 133932 78752 133938 78804
rect 135990 78752 135996 78804
rect 136048 78792 136054 78804
rect 136174 78792 136180 78804
rect 136048 78764 136180 78792
rect 136048 78752 136054 78764
rect 136174 78752 136180 78764
rect 136232 78752 136238 78804
rect 140746 78792 140774 78832
rect 154206 78820 154212 78832
rect 154264 78820 154270 78872
rect 136284 78764 138014 78792
rect 140746 78764 149054 78792
rect 130838 78684 130844 78736
rect 130896 78724 130902 78736
rect 136284 78724 136312 78764
rect 130896 78696 136312 78724
rect 130896 78684 130902 78696
rect 122156 78628 125594 78656
rect 137986 78656 138014 78764
rect 138566 78684 138572 78736
rect 138624 78724 138630 78736
rect 139210 78724 139216 78736
rect 138624 78696 139216 78724
rect 138624 78684 138630 78696
rect 139210 78684 139216 78696
rect 139268 78684 139274 78736
rect 140038 78684 140044 78736
rect 140096 78724 140102 78736
rect 140498 78724 140504 78736
rect 140096 78696 140504 78724
rect 140096 78684 140102 78696
rect 140498 78684 140504 78696
rect 140556 78684 140562 78736
rect 144362 78656 144368 78668
rect 137986 78628 144368 78656
rect 122156 78616 122162 78628
rect 144362 78616 144368 78628
rect 144420 78616 144426 78668
rect 149026 78656 149054 78764
rect 155218 78684 155224 78736
rect 155276 78724 155282 78736
rect 155328 78724 155356 78888
rect 158806 78820 158812 78872
rect 158864 78860 158870 78872
rect 170232 78860 170260 78900
rect 158864 78832 170260 78860
rect 171750 78860 171778 78900
rect 172882 78888 172888 78940
rect 172940 78928 172946 78940
rect 173158 78928 173164 78940
rect 172940 78900 173164 78928
rect 172940 78888 172946 78900
rect 173158 78888 173164 78900
rect 173216 78888 173222 78940
rect 174464 78928 174492 78968
rect 176194 78956 176200 79008
rect 176252 78996 176258 79008
rect 192754 78996 192760 79008
rect 176252 78968 192760 78996
rect 176252 78956 176258 78968
rect 192754 78956 192760 78968
rect 192812 78956 192818 79008
rect 178586 78928 178592 78940
rect 174464 78900 178592 78928
rect 178586 78888 178592 78900
rect 178644 78888 178650 78940
rect 177850 78860 177856 78872
rect 171750 78832 177856 78860
rect 158864 78820 158870 78832
rect 177850 78820 177856 78832
rect 177908 78820 177914 78872
rect 178034 78820 178040 78872
rect 178092 78860 178098 78872
rect 180518 78860 180524 78872
rect 178092 78832 180524 78860
rect 178092 78820 178098 78832
rect 180518 78820 180524 78832
rect 180576 78820 180582 78872
rect 158530 78792 158536 78804
rect 155276 78696 155356 78724
rect 156616 78764 158536 78792
rect 155276 78684 155282 78696
rect 156616 78656 156644 78764
rect 158530 78752 158536 78764
rect 158588 78752 158594 78804
rect 162394 78752 162400 78804
rect 162452 78792 162458 78804
rect 162452 78764 162716 78792
rect 162452 78752 162458 78764
rect 162688 78736 162716 78764
rect 164786 78752 164792 78804
rect 164844 78792 164850 78804
rect 169570 78792 169576 78804
rect 164844 78764 169576 78792
rect 164844 78752 164850 78764
rect 169570 78752 169576 78764
rect 169628 78752 169634 78804
rect 170122 78752 170128 78804
rect 170180 78792 170186 78804
rect 178402 78792 178408 78804
rect 170180 78764 178408 78792
rect 170180 78752 170186 78764
rect 178402 78752 178408 78764
rect 178460 78752 178466 78804
rect 157334 78684 157340 78736
rect 157392 78724 157398 78736
rect 161106 78724 161112 78736
rect 157392 78696 161112 78724
rect 157392 78684 157398 78696
rect 161106 78684 161112 78696
rect 161164 78684 161170 78736
rect 161198 78684 161204 78736
rect 161256 78724 161262 78736
rect 162578 78724 162584 78736
rect 161256 78696 162584 78724
rect 161256 78684 161262 78696
rect 162578 78684 162584 78696
rect 162636 78684 162642 78736
rect 162670 78684 162676 78736
rect 162728 78684 162734 78736
rect 167178 78684 167184 78736
rect 167236 78724 167242 78736
rect 167454 78724 167460 78736
rect 167236 78696 167460 78724
rect 167236 78684 167242 78696
rect 167454 78684 167460 78696
rect 167512 78684 167518 78736
rect 177758 78724 177764 78736
rect 170600 78696 177764 78724
rect 149026 78628 156644 78656
rect 161014 78616 161020 78668
rect 161072 78656 161078 78668
rect 162394 78656 162400 78668
rect 161072 78628 162400 78656
rect 161072 78616 161078 78628
rect 162394 78616 162400 78628
rect 162452 78616 162458 78668
rect 164234 78616 164240 78668
rect 164292 78656 164298 78668
rect 164418 78656 164424 78668
rect 164292 78628 164424 78656
rect 164292 78616 164298 78628
rect 164418 78616 164424 78628
rect 164476 78616 164482 78668
rect 164602 78616 164608 78668
rect 164660 78656 164666 78668
rect 164786 78656 164792 78668
rect 164660 78628 164792 78656
rect 164660 78616 164666 78628
rect 164786 78616 164792 78628
rect 164844 78616 164850 78668
rect 166166 78616 166172 78668
rect 166224 78656 166230 78668
rect 170122 78656 170128 78668
rect 166224 78628 170128 78656
rect 166224 78616 166230 78628
rect 170122 78616 170128 78628
rect 170180 78616 170186 78668
rect 150710 78548 150716 78600
rect 150768 78588 150774 78600
rect 170600 78588 170628 78696
rect 177758 78684 177764 78696
rect 177816 78684 177822 78736
rect 171594 78616 171600 78668
rect 171652 78656 171658 78668
rect 174814 78656 174820 78668
rect 171652 78628 174820 78656
rect 171652 78616 171658 78628
rect 174814 78616 174820 78628
rect 174872 78616 174878 78668
rect 175826 78616 175832 78668
rect 175884 78656 175890 78668
rect 177206 78656 177212 78668
rect 175884 78628 177212 78656
rect 175884 78616 175890 78628
rect 177206 78616 177212 78628
rect 177264 78616 177270 78668
rect 177390 78616 177396 78668
rect 177448 78656 177454 78668
rect 177448 78628 183554 78656
rect 177448 78616 177454 78628
rect 150768 78560 170628 78588
rect 150768 78548 150774 78560
rect 173066 78548 173072 78600
rect 173124 78588 173130 78600
rect 178770 78588 178776 78600
rect 173124 78560 178776 78588
rect 173124 78548 173130 78560
rect 178770 78548 178776 78560
rect 178828 78548 178834 78600
rect 183526 78588 183554 78628
rect 580626 78588 580632 78600
rect 183526 78560 580632 78588
rect 580626 78548 580632 78560
rect 580684 78548 580690 78600
rect 134426 78480 134432 78532
rect 134484 78520 134490 78532
rect 134794 78520 134800 78532
rect 134484 78492 134800 78520
rect 134484 78480 134490 78492
rect 134794 78480 134800 78492
rect 134852 78480 134858 78532
rect 136358 78480 136364 78532
rect 136416 78520 136422 78532
rect 137186 78520 137192 78532
rect 136416 78492 137192 78520
rect 136416 78480 136422 78492
rect 137186 78480 137192 78492
rect 137244 78480 137250 78532
rect 146570 78480 146576 78532
rect 146628 78520 146634 78532
rect 171042 78520 171048 78532
rect 146628 78492 171048 78520
rect 146628 78480 146634 78492
rect 171042 78480 171048 78492
rect 171100 78480 171106 78532
rect 172882 78480 172888 78532
rect 172940 78520 172946 78532
rect 173802 78520 173808 78532
rect 172940 78492 173808 78520
rect 172940 78480 172946 78492
rect 173802 78480 173808 78492
rect 173860 78480 173866 78532
rect 175642 78480 175648 78532
rect 175700 78520 175706 78532
rect 176562 78520 176568 78532
rect 175700 78492 176568 78520
rect 175700 78480 175706 78492
rect 176562 78480 176568 78492
rect 176620 78480 176626 78532
rect 176746 78480 176752 78532
rect 176804 78520 176810 78532
rect 179138 78520 179144 78532
rect 176804 78492 179144 78520
rect 176804 78480 176810 78492
rect 179138 78480 179144 78492
rect 179196 78480 179202 78532
rect 180242 78480 180248 78532
rect 180300 78520 180306 78532
rect 188890 78520 188896 78532
rect 180300 78492 188896 78520
rect 180300 78480 180306 78492
rect 188890 78480 188896 78492
rect 188948 78480 188954 78532
rect 130654 78412 130660 78464
rect 130712 78452 130718 78464
rect 138658 78452 138664 78464
rect 130712 78424 138664 78452
rect 130712 78412 130718 78424
rect 138658 78412 138664 78424
rect 138716 78412 138722 78464
rect 140130 78412 140136 78464
rect 140188 78452 140194 78464
rect 154574 78452 154580 78464
rect 140188 78424 154580 78452
rect 140188 78412 140194 78424
rect 154574 78412 154580 78424
rect 154632 78412 154638 78464
rect 161566 78412 161572 78464
rect 161624 78452 161630 78464
rect 162026 78452 162032 78464
rect 161624 78424 162032 78452
rect 161624 78412 161630 78424
rect 162026 78412 162032 78424
rect 162084 78412 162090 78464
rect 164050 78412 164056 78464
rect 164108 78452 164114 78464
rect 171502 78452 171508 78464
rect 164108 78424 171508 78452
rect 164108 78412 164114 78424
rect 171502 78412 171508 78424
rect 171560 78412 171566 78464
rect 454034 78452 454040 78464
rect 171612 78424 454040 78452
rect 158714 78344 158720 78396
rect 158772 78384 158778 78396
rect 163958 78384 163964 78396
rect 158772 78356 163964 78384
rect 158772 78344 158778 78356
rect 163958 78344 163964 78356
rect 164016 78344 164022 78396
rect 170122 78344 170128 78396
rect 170180 78384 170186 78396
rect 171612 78384 171640 78424
rect 454034 78412 454040 78424
rect 454092 78412 454098 78464
rect 170180 78356 171640 78384
rect 170180 78344 170186 78356
rect 171778 78344 171784 78396
rect 171836 78384 171842 78396
rect 460934 78384 460940 78396
rect 171836 78356 460940 78384
rect 171836 78344 171842 78356
rect 460934 78344 460940 78356
rect 460992 78344 460998 78396
rect 129458 78276 129464 78328
rect 129516 78316 129522 78328
rect 139578 78316 139584 78328
rect 129516 78288 139584 78316
rect 129516 78276 129522 78288
rect 139578 78276 139584 78288
rect 139636 78276 139642 78328
rect 140130 78276 140136 78328
rect 140188 78316 140194 78328
rect 140866 78316 140872 78328
rect 140188 78288 140872 78316
rect 140188 78276 140194 78288
rect 140866 78276 140872 78288
rect 140924 78276 140930 78328
rect 161382 78276 161388 78328
rect 161440 78316 161446 78328
rect 166166 78316 166172 78328
rect 161440 78288 166172 78316
rect 161440 78276 161446 78288
rect 166166 78276 166172 78288
rect 166224 78276 166230 78328
rect 167362 78276 167368 78328
rect 167420 78316 167426 78328
rect 467834 78316 467840 78328
rect 167420 78288 467840 78316
rect 167420 78276 167426 78288
rect 467834 78276 467840 78288
rect 467892 78276 467898 78328
rect 127710 78208 127716 78260
rect 127768 78248 127774 78260
rect 134518 78248 134524 78260
rect 127768 78220 134524 78248
rect 127768 78208 127774 78220
rect 134518 78208 134524 78220
rect 134576 78208 134582 78260
rect 161658 78208 161664 78260
rect 161716 78248 161722 78260
rect 162670 78248 162676 78260
rect 161716 78220 162676 78248
rect 161716 78208 161722 78220
rect 162670 78208 162676 78220
rect 162728 78208 162734 78260
rect 167546 78208 167552 78260
rect 167604 78248 167610 78260
rect 474734 78248 474740 78260
rect 167604 78220 474740 78248
rect 167604 78208 167610 78220
rect 474734 78208 474740 78220
rect 474792 78208 474798 78260
rect 118694 78140 118700 78192
rect 118752 78180 118758 78192
rect 139394 78180 139400 78192
rect 118752 78152 139400 78180
rect 118752 78140 118758 78152
rect 139394 78140 139400 78152
rect 139452 78140 139458 78192
rect 157794 78140 157800 78192
rect 157852 78180 157858 78192
rect 164602 78180 164608 78192
rect 157852 78152 164608 78180
rect 157852 78140 157858 78152
rect 164602 78140 164608 78152
rect 164660 78140 164666 78192
rect 172606 78140 172612 78192
rect 172664 78180 172670 78192
rect 172974 78180 172980 78192
rect 172664 78152 172980 78180
rect 172664 78140 172670 78152
rect 172974 78140 172980 78152
rect 173032 78140 173038 78192
rect 175366 78140 175372 78192
rect 175424 78180 175430 78192
rect 175424 78152 179736 78180
rect 175424 78140 175430 78152
rect 96614 78072 96620 78124
rect 96672 78112 96678 78124
rect 138014 78112 138020 78124
rect 96672 78084 138020 78112
rect 96672 78072 96678 78084
rect 138014 78072 138020 78084
rect 138072 78072 138078 78124
rect 145466 78072 145472 78124
rect 145524 78112 145530 78124
rect 147306 78112 147312 78124
rect 145524 78084 147312 78112
rect 145524 78072 145530 78084
rect 147306 78072 147312 78084
rect 147364 78072 147370 78124
rect 150802 78072 150808 78124
rect 150860 78112 150866 78124
rect 150860 78084 158714 78112
rect 150860 78072 150866 78084
rect 78674 78004 78680 78056
rect 78732 78044 78738 78056
rect 136818 78044 136824 78056
rect 78732 78016 136824 78044
rect 78732 78004 78738 78016
rect 136818 78004 136824 78016
rect 136876 78004 136882 78056
rect 145190 78004 145196 78056
rect 145248 78044 145254 78056
rect 158686 78044 158714 78084
rect 159910 78072 159916 78124
rect 159968 78112 159974 78124
rect 165798 78112 165804 78124
rect 159968 78084 165804 78112
rect 159968 78072 159974 78084
rect 165798 78072 165804 78084
rect 165856 78072 165862 78124
rect 170306 78072 170312 78124
rect 170364 78112 170370 78124
rect 170364 78084 175688 78112
rect 170364 78072 170370 78084
rect 145248 78016 151814 78044
rect 158686 78016 162164 78044
rect 145248 78004 145254 78016
rect 10318 77936 10324 77988
rect 10376 77976 10382 77988
rect 129550 77976 129556 77988
rect 10376 77948 129556 77976
rect 10376 77936 10382 77948
rect 129550 77936 129556 77948
rect 129608 77936 129614 77988
rect 131482 77936 131488 77988
rect 131540 77976 131546 77988
rect 132402 77976 132408 77988
rect 131540 77948 132408 77976
rect 131540 77936 131546 77948
rect 132402 77936 132408 77948
rect 132460 77936 132466 77988
rect 145374 77936 145380 77988
rect 145432 77976 145438 77988
rect 147582 77976 147588 77988
rect 145432 77948 147588 77976
rect 145432 77936 145438 77948
rect 147582 77936 147588 77948
rect 147640 77936 147646 77988
rect 151786 77976 151814 78016
rect 151786 77948 161106 77976
rect 131666 77868 131672 77920
rect 131724 77908 131730 77920
rect 131942 77908 131948 77920
rect 131724 77880 131948 77908
rect 131724 77868 131730 77880
rect 131942 77868 131948 77880
rect 132000 77868 132006 77920
rect 128998 77800 129004 77852
rect 129056 77840 129062 77852
rect 135254 77840 135260 77852
rect 129056 77812 135260 77840
rect 129056 77800 129062 77812
rect 135254 77800 135260 77812
rect 135312 77800 135318 77852
rect 129182 77732 129188 77784
rect 129240 77772 129246 77784
rect 139026 77772 139032 77784
rect 129240 77744 139032 77772
rect 129240 77732 129246 77744
rect 139026 77732 139032 77744
rect 139084 77732 139090 77784
rect 128354 77664 128360 77716
rect 128412 77704 128418 77716
rect 140774 77704 140780 77716
rect 128412 77676 140780 77704
rect 128412 77664 128418 77676
rect 140774 77664 140780 77676
rect 140832 77664 140838 77716
rect 161078 77704 161106 77948
rect 162136 77840 162164 78016
rect 172698 78004 172704 78056
rect 172756 78044 172762 78056
rect 172974 78044 172980 78056
rect 172756 78016 172980 78044
rect 172756 78004 172762 78016
rect 172974 78004 172980 78016
rect 173032 78004 173038 78056
rect 173986 78004 173992 78056
rect 174044 78044 174050 78056
rect 174446 78044 174452 78056
rect 174044 78016 174452 78044
rect 174044 78004 174050 78016
rect 174446 78004 174452 78016
rect 174504 78004 174510 78056
rect 175660 78044 175688 78084
rect 175734 78072 175740 78124
rect 175792 78112 175798 78124
rect 179708 78112 179736 78152
rect 179874 78140 179880 78192
rect 179932 78180 179938 78192
rect 557534 78180 557540 78192
rect 179932 78152 557540 78180
rect 179932 78140 179938 78152
rect 557534 78140 557540 78152
rect 557592 78140 557598 78192
rect 574094 78112 574100 78124
rect 175792 78084 179644 78112
rect 179708 78084 574100 78112
rect 175792 78072 175798 78084
rect 175826 78044 175832 78056
rect 175660 78016 175832 78044
rect 175826 78004 175832 78016
rect 175884 78004 175890 78056
rect 179616 78044 179644 78084
rect 574094 78072 574100 78084
rect 574152 78072 574158 78124
rect 580994 78044 581000 78056
rect 179616 78016 581000 78044
rect 580994 78004 581000 78016
rect 581052 78004 581058 78056
rect 162854 77936 162860 77988
rect 162912 77976 162918 77988
rect 162912 77948 171548 77976
rect 162912 77936 162918 77948
rect 162210 77868 162216 77920
rect 162268 77908 162274 77920
rect 171520 77908 171548 77948
rect 173434 77936 173440 77988
rect 173492 77976 173498 77988
rect 175918 77976 175924 77988
rect 173492 77948 175924 77976
rect 173492 77936 173498 77948
rect 175918 77936 175924 77948
rect 175976 77936 175982 77988
rect 176470 77936 176476 77988
rect 176528 77976 176534 77988
rect 187878 77976 187884 77988
rect 176528 77948 187884 77976
rect 176528 77936 176534 77948
rect 187878 77936 187884 77948
rect 187936 77936 187942 77988
rect 582374 77976 582380 77988
rect 191024 77948 582380 77976
rect 176194 77908 176200 77920
rect 162268 77880 171456 77908
rect 171520 77880 176200 77908
rect 162268 77868 162274 77880
rect 162136 77812 166994 77840
rect 166966 77772 166994 77812
rect 168190 77772 168196 77784
rect 166966 77744 168196 77772
rect 168190 77732 168196 77744
rect 168248 77732 168254 77784
rect 171428 77772 171456 77880
rect 176194 77868 176200 77880
rect 176252 77868 176258 77920
rect 177206 77868 177212 77920
rect 177264 77908 177270 77920
rect 191024 77908 191052 77948
rect 582374 77936 582380 77948
rect 582432 77936 582438 77988
rect 580166 77908 580172 77920
rect 177264 77880 191052 77908
rect 193186 77880 580172 77908
rect 177264 77868 177270 77880
rect 171502 77800 171508 77852
rect 171560 77840 171566 77852
rect 177298 77840 177304 77852
rect 171560 77812 177304 77840
rect 171560 77800 171566 77812
rect 177298 77800 177304 77812
rect 177356 77800 177362 77852
rect 187878 77800 187884 77852
rect 187936 77840 187942 77852
rect 193186 77840 193214 77880
rect 580166 77868 580172 77880
rect 580224 77868 580230 77920
rect 187936 77812 193214 77840
rect 187936 77800 187942 77812
rect 176378 77772 176384 77784
rect 171428 77744 176384 77772
rect 176378 77732 176384 77744
rect 176436 77732 176442 77784
rect 161078 77676 166994 77704
rect 129826 77596 129832 77648
rect 129884 77636 129890 77648
rect 136726 77636 136732 77648
rect 129884 77608 136732 77636
rect 129884 77596 129890 77608
rect 136726 77596 136732 77608
rect 136784 77596 136790 77648
rect 148042 77596 148048 77648
rect 148100 77636 148106 77648
rect 148410 77636 148416 77648
rect 148100 77608 148416 77636
rect 148100 77596 148106 77608
rect 148410 77596 148416 77608
rect 148468 77596 148474 77648
rect 166966 77636 166994 77676
rect 169570 77664 169576 77716
rect 169628 77704 169634 77716
rect 177206 77704 177212 77716
rect 169628 77676 177212 77704
rect 169628 77664 169634 77676
rect 177206 77664 177212 77676
rect 177264 77664 177270 77716
rect 172422 77636 172428 77648
rect 166966 77608 172428 77636
rect 172422 77596 172428 77608
rect 172480 77596 172486 77648
rect 174814 77596 174820 77648
rect 174872 77636 174878 77648
rect 178770 77636 178776 77648
rect 174872 77608 178776 77636
rect 174872 77596 174878 77608
rect 178770 77596 178776 77608
rect 178828 77596 178834 77648
rect 130746 77528 130752 77580
rect 130804 77568 130810 77580
rect 132126 77568 132132 77580
rect 130804 77540 132132 77568
rect 130804 77528 130810 77540
rect 132126 77528 132132 77540
rect 132184 77528 132190 77580
rect 135254 77528 135260 77580
rect 135312 77568 135318 77580
rect 140866 77568 140872 77580
rect 135312 77540 140872 77568
rect 135312 77528 135318 77540
rect 140866 77528 140872 77540
rect 140924 77528 140930 77580
rect 147950 77528 147956 77580
rect 148008 77568 148014 77580
rect 148226 77568 148232 77580
rect 148008 77540 148232 77568
rect 148008 77528 148014 77540
rect 148226 77528 148232 77540
rect 148284 77528 148290 77580
rect 148686 77528 148692 77580
rect 148744 77568 148750 77580
rect 172330 77568 172336 77580
rect 148744 77540 172336 77568
rect 148744 77528 148750 77540
rect 172330 77528 172336 77540
rect 172388 77528 172394 77580
rect 180610 77528 180616 77580
rect 180668 77568 180674 77580
rect 190454 77568 190460 77580
rect 180668 77540 190460 77568
rect 180668 77528 180674 77540
rect 190454 77528 190460 77540
rect 190512 77528 190518 77580
rect 131850 77460 131856 77512
rect 131908 77500 131914 77512
rect 135622 77500 135628 77512
rect 131908 77472 135628 77500
rect 131908 77460 131914 77472
rect 135622 77460 135628 77472
rect 135680 77460 135686 77512
rect 156138 77460 156144 77512
rect 156196 77500 156202 77512
rect 168282 77500 168288 77512
rect 156196 77472 168288 77500
rect 156196 77460 156202 77472
rect 168282 77460 168288 77472
rect 168340 77460 168346 77512
rect 171042 77460 171048 77512
rect 171100 77500 171106 77512
rect 177482 77500 177488 77512
rect 171100 77472 177488 77500
rect 171100 77460 171106 77472
rect 177482 77460 177488 77472
rect 177540 77460 177546 77512
rect 129274 77392 129280 77444
rect 129332 77432 129338 77444
rect 132034 77432 132040 77444
rect 129332 77404 132040 77432
rect 129332 77392 129338 77404
rect 132034 77392 132040 77404
rect 132092 77392 132098 77444
rect 132126 77392 132132 77444
rect 132184 77432 132190 77444
rect 133138 77432 133144 77444
rect 132184 77404 133144 77432
rect 132184 77392 132190 77404
rect 133138 77392 133144 77404
rect 133196 77392 133202 77444
rect 140682 77392 140688 77444
rect 140740 77432 140746 77444
rect 143166 77432 143172 77444
rect 140740 77404 143172 77432
rect 140740 77392 140746 77404
rect 143166 77392 143172 77404
rect 143224 77392 143230 77444
rect 143718 77392 143724 77444
rect 143776 77432 143782 77444
rect 144362 77432 144368 77444
rect 143776 77404 144368 77432
rect 143776 77392 143782 77404
rect 144362 77392 144368 77404
rect 144420 77392 144426 77444
rect 157886 77392 157892 77444
rect 157944 77432 157950 77444
rect 158806 77432 158812 77444
rect 157944 77404 158812 77432
rect 157944 77392 157950 77404
rect 158806 77392 158812 77404
rect 158864 77392 158870 77444
rect 160370 77392 160376 77444
rect 160428 77432 160434 77444
rect 165430 77432 165436 77444
rect 160428 77404 165436 77432
rect 160428 77392 160434 77404
rect 165430 77392 165436 77404
rect 165488 77392 165494 77444
rect 168374 77392 168380 77444
rect 168432 77432 168438 77444
rect 173802 77432 173808 77444
rect 168432 77404 173808 77432
rect 168432 77392 168438 77404
rect 173802 77392 173808 77404
rect 173860 77392 173866 77444
rect 130378 77324 130384 77376
rect 130436 77364 130442 77376
rect 137830 77364 137836 77376
rect 130436 77336 137836 77364
rect 130436 77324 130442 77336
rect 137830 77324 137836 77336
rect 137888 77324 137894 77376
rect 164326 77324 164332 77376
rect 164384 77364 164390 77376
rect 177666 77364 177672 77376
rect 164384 77336 177672 77364
rect 164384 77324 164390 77336
rect 177666 77324 177672 77336
rect 177724 77324 177730 77376
rect 126238 77256 126244 77308
rect 126296 77296 126302 77308
rect 130562 77296 130568 77308
rect 126296 77268 130568 77296
rect 126296 77256 126302 77268
rect 130562 77256 130568 77268
rect 130620 77256 130626 77308
rect 132402 77256 132408 77308
rect 132460 77296 132466 77308
rect 134242 77296 134248 77308
rect 132460 77268 134248 77296
rect 132460 77256 132466 77268
rect 134242 77256 134248 77268
rect 134300 77256 134306 77308
rect 134518 77256 134524 77308
rect 134576 77296 134582 77308
rect 136450 77296 136456 77308
rect 134576 77268 136456 77296
rect 134576 77256 134582 77268
rect 136450 77256 136456 77268
rect 136508 77256 136514 77308
rect 163682 77256 163688 77308
rect 163740 77296 163746 77308
rect 165338 77296 165344 77308
rect 163740 77268 165344 77296
rect 163740 77256 163746 77268
rect 165338 77256 165344 77268
rect 165396 77256 165402 77308
rect 165798 77256 165804 77308
rect 165856 77296 165862 77308
rect 166626 77296 166632 77308
rect 165856 77268 166632 77296
rect 165856 77256 165862 77268
rect 166626 77256 166632 77268
rect 166684 77256 166690 77308
rect 178218 77256 178224 77308
rect 178276 77296 178282 77308
rect 179782 77296 179788 77308
rect 178276 77268 179788 77296
rect 178276 77256 178282 77268
rect 179782 77256 179788 77268
rect 179840 77256 179846 77308
rect 126974 77188 126980 77240
rect 127032 77228 127038 77240
rect 140406 77228 140412 77240
rect 127032 77200 140412 77228
rect 127032 77188 127038 77200
rect 140406 77188 140412 77200
rect 140464 77188 140470 77240
rect 144822 77188 144828 77240
rect 144880 77228 144886 77240
rect 185026 77228 185032 77240
rect 144880 77200 185032 77228
rect 144880 77188 144886 77200
rect 185026 77188 185032 77200
rect 185084 77188 185090 77240
rect 132420 77132 137784 77160
rect 104894 76984 104900 77036
rect 104952 77024 104958 77036
rect 132420 77024 132448 77132
rect 104952 76996 132448 77024
rect 137756 77024 137784 77132
rect 145098 77120 145104 77172
rect 145156 77160 145162 77172
rect 145742 77160 145748 77172
rect 145156 77132 145748 77160
rect 145156 77120 145162 77132
rect 145742 77120 145748 77132
rect 145800 77120 145806 77172
rect 146202 77120 146208 77172
rect 146260 77160 146266 77172
rect 147674 77160 147680 77172
rect 146260 77132 147680 77160
rect 146260 77120 146266 77132
rect 147674 77120 147680 77132
rect 147732 77120 147738 77172
rect 147766 77120 147772 77172
rect 147824 77160 147830 77172
rect 148042 77160 148048 77172
rect 147824 77132 148048 77160
rect 147824 77120 147830 77132
rect 148042 77120 148048 77132
rect 148100 77120 148106 77172
rect 173066 77120 173072 77172
rect 173124 77160 173130 77172
rect 173618 77160 173624 77172
rect 173124 77132 173624 77160
rect 173124 77120 173130 77132
rect 173618 77120 173624 77132
rect 173676 77120 173682 77172
rect 175274 77120 175280 77172
rect 175332 77160 175338 77172
rect 233234 77160 233240 77172
rect 175332 77132 233240 77160
rect 175332 77120 175338 77132
rect 233234 77120 233240 77132
rect 233292 77120 233298 77172
rect 155402 77052 155408 77104
rect 155460 77092 155466 77104
rect 222930 77092 222936 77104
rect 155460 77064 222936 77092
rect 155460 77052 155466 77064
rect 222930 77052 222936 77064
rect 222988 77052 222994 77104
rect 138842 77024 138848 77036
rect 137756 76996 138848 77024
rect 104952 76984 104958 76996
rect 138842 76984 138848 76996
rect 138900 76984 138906 77036
rect 150618 76984 150624 77036
rect 150676 77024 150682 77036
rect 150894 77024 150900 77036
rect 150676 76996 150900 77024
rect 150676 76984 150682 76996
rect 150894 76984 150900 76996
rect 150952 76984 150958 77036
rect 168190 76984 168196 77036
rect 168248 77024 168254 77036
rect 259454 77024 259460 77036
rect 168248 76996 259460 77024
rect 168248 76984 168254 76996
rect 259454 76984 259460 76996
rect 259512 76984 259518 77036
rect 91094 76916 91100 76968
rect 91152 76956 91158 76968
rect 137646 76956 137652 76968
rect 91152 76928 137652 76956
rect 91152 76916 91158 76928
rect 137646 76916 137652 76928
rect 137704 76916 137710 76968
rect 145374 76916 145380 76968
rect 145432 76956 145438 76968
rect 146110 76956 146116 76968
rect 145432 76928 146116 76956
rect 145432 76916 145438 76928
rect 146110 76916 146116 76928
rect 146168 76916 146174 76968
rect 153286 76916 153292 76968
rect 153344 76956 153350 76968
rect 153746 76956 153752 76968
rect 153344 76928 153752 76956
rect 153344 76916 153350 76928
rect 153746 76916 153752 76928
rect 153804 76916 153810 76968
rect 159358 76916 159364 76968
rect 159416 76956 159422 76968
rect 273530 76956 273536 76968
rect 159416 76928 273536 76956
rect 159416 76916 159422 76928
rect 273530 76916 273536 76928
rect 273588 76916 273594 76968
rect 85574 76848 85580 76900
rect 85632 76888 85638 76900
rect 136358 76888 136364 76900
rect 85632 76860 136364 76888
rect 85632 76848 85638 76860
rect 136358 76848 136364 76860
rect 136416 76848 136422 76900
rect 151446 76848 151452 76900
rect 151504 76888 151510 76900
rect 267734 76888 267740 76900
rect 151504 76860 267740 76888
rect 151504 76848 151510 76860
rect 267734 76848 267740 76860
rect 267792 76848 267798 76900
rect 84194 76780 84200 76832
rect 84252 76820 84258 76832
rect 136634 76820 136640 76832
rect 84252 76792 136640 76820
rect 84252 76780 84258 76792
rect 136634 76780 136640 76792
rect 136692 76780 136698 76832
rect 160278 76780 160284 76832
rect 160336 76820 160342 76832
rect 280338 76820 280344 76832
rect 160336 76792 280344 76820
rect 160336 76780 160342 76792
rect 280338 76780 280344 76792
rect 280396 76780 280402 76832
rect 67634 76712 67640 76764
rect 67692 76752 67698 76764
rect 131850 76752 131856 76764
rect 67692 76724 131856 76752
rect 67692 76712 67698 76724
rect 131850 76712 131856 76724
rect 131908 76712 131914 76764
rect 142338 76712 142344 76764
rect 142396 76752 142402 76764
rect 143074 76752 143080 76764
rect 142396 76724 143080 76752
rect 142396 76712 142402 76724
rect 143074 76712 143080 76724
rect 143132 76712 143138 76764
rect 160646 76712 160652 76764
rect 160704 76752 160710 76764
rect 311894 76752 311900 76764
rect 160704 76724 311900 76752
rect 160704 76712 160710 76724
rect 311894 76712 311900 76724
rect 311952 76712 311958 76764
rect 59354 76644 59360 76696
rect 59412 76684 59418 76696
rect 135162 76684 135168 76696
rect 59412 76656 135168 76684
rect 59412 76644 59418 76656
rect 135162 76644 135168 76656
rect 135220 76644 135226 76696
rect 158898 76644 158904 76696
rect 158956 76684 158962 76696
rect 336734 76684 336740 76696
rect 158956 76656 336740 76684
rect 158956 76644 158962 76656
rect 336734 76644 336740 76656
rect 336792 76644 336798 76696
rect 34514 76576 34520 76628
rect 34572 76616 34578 76628
rect 34572 76588 129734 76616
rect 34572 76576 34578 76588
rect 11054 76508 11060 76560
rect 11112 76548 11118 76560
rect 127158 76548 127164 76560
rect 11112 76520 127164 76548
rect 11112 76508 11118 76520
rect 127158 76508 127164 76520
rect 127216 76508 127222 76560
rect 129706 76480 129734 76588
rect 133046 76576 133052 76628
rect 133104 76616 133110 76628
rect 133506 76616 133512 76628
rect 133104 76588 133512 76616
rect 133104 76576 133110 76588
rect 133506 76576 133512 76588
rect 133564 76576 133570 76628
rect 142154 76576 142160 76628
rect 142212 76616 142218 76628
rect 142614 76616 142620 76628
rect 142212 76588 142620 76616
rect 142212 76576 142218 76588
rect 142614 76576 142620 76588
rect 142672 76576 142678 76628
rect 142706 76576 142712 76628
rect 142764 76616 142770 76628
rect 142890 76616 142896 76628
rect 142764 76588 142896 76616
rect 142764 76576 142770 76588
rect 142890 76576 142896 76588
rect 142948 76576 142954 76628
rect 147674 76576 147680 76628
rect 147732 76616 147738 76628
rect 148502 76616 148508 76628
rect 147732 76588 148508 76616
rect 147732 76576 147738 76588
rect 148502 76576 148508 76588
rect 148560 76576 148566 76628
rect 160278 76576 160284 76628
rect 160336 76616 160342 76628
rect 160738 76616 160744 76628
rect 160336 76588 160744 76616
rect 160336 76576 160342 76588
rect 160738 76576 160744 76588
rect 160796 76576 160802 76628
rect 172790 76576 172796 76628
rect 172848 76616 172854 76628
rect 173158 76616 173164 76628
rect 172848 76588 173164 76616
rect 172848 76576 172854 76588
rect 173158 76576 173164 76588
rect 173216 76576 173222 76628
rect 177850 76576 177856 76628
rect 177908 76616 177914 76628
rect 361574 76616 361580 76628
rect 177908 76588 361580 76616
rect 177908 76576 177914 76588
rect 361574 76576 361580 76588
rect 361632 76576 361638 76628
rect 132678 76508 132684 76560
rect 132736 76548 132742 76560
rect 133690 76548 133696 76560
rect 132736 76520 133696 76548
rect 132736 76508 132742 76520
rect 133690 76508 133696 76520
rect 133748 76508 133754 76560
rect 147122 76508 147128 76560
rect 147180 76548 147186 76560
rect 148134 76548 148140 76560
rect 147180 76520 148140 76548
rect 147180 76508 147186 76520
rect 148134 76508 148140 76520
rect 148192 76508 148198 76560
rect 149606 76508 149612 76560
rect 149664 76548 149670 76560
rect 150066 76548 150072 76560
rect 149664 76520 150072 76548
rect 149664 76508 149670 76520
rect 150066 76508 150072 76520
rect 150124 76508 150130 76560
rect 161842 76508 161848 76560
rect 161900 76548 161906 76560
rect 398834 76548 398840 76560
rect 161900 76520 398840 76548
rect 161900 76508 161906 76520
rect 398834 76508 398840 76520
rect 398892 76508 398898 76560
rect 133230 76480 133236 76492
rect 129706 76452 133236 76480
rect 133230 76440 133236 76452
rect 133288 76440 133294 76492
rect 156690 76440 156696 76492
rect 156748 76480 156754 76492
rect 178494 76480 178500 76492
rect 156748 76452 178500 76480
rect 156748 76440 156754 76452
rect 178494 76440 178500 76452
rect 178552 76440 178558 76492
rect 131482 76372 131488 76424
rect 131540 76412 131546 76424
rect 132218 76412 132224 76424
rect 131540 76384 132224 76412
rect 131540 76372 131546 76384
rect 132218 76372 132224 76384
rect 132276 76372 132282 76424
rect 145466 76372 145472 76424
rect 145524 76412 145530 76424
rect 146018 76412 146024 76424
rect 145524 76384 146024 76412
rect 145524 76372 145530 76384
rect 146018 76372 146024 76384
rect 146076 76372 146082 76424
rect 149606 76372 149612 76424
rect 149664 76412 149670 76424
rect 149882 76412 149888 76424
rect 149664 76384 149888 76412
rect 149664 76372 149670 76384
rect 149882 76372 149888 76384
rect 149940 76372 149946 76424
rect 156414 76372 156420 76424
rect 156472 76412 156478 76424
rect 156472 76384 171824 76412
rect 156472 76372 156478 76384
rect 143810 76304 143816 76356
rect 143868 76344 143874 76356
rect 144086 76344 144092 76356
rect 143868 76316 144092 76344
rect 143868 76304 143874 76316
rect 144086 76304 144092 76316
rect 144144 76304 144150 76356
rect 164602 76304 164608 76356
rect 164660 76344 164666 76356
rect 165246 76344 165252 76356
rect 164660 76316 165252 76344
rect 164660 76304 164666 76316
rect 165246 76304 165252 76316
rect 165304 76304 165310 76356
rect 146386 76236 146392 76288
rect 146444 76276 146450 76288
rect 149882 76276 149888 76288
rect 146444 76248 149888 76276
rect 146444 76236 146450 76248
rect 149882 76236 149888 76248
rect 149940 76236 149946 76288
rect 153378 76236 153384 76288
rect 153436 76276 153442 76288
rect 153562 76276 153568 76288
rect 153436 76248 153568 76276
rect 153436 76236 153442 76248
rect 153562 76236 153568 76248
rect 153620 76236 153626 76288
rect 169846 76236 169852 76288
rect 169904 76276 169910 76288
rect 170306 76276 170312 76288
rect 169904 76248 170312 76276
rect 169904 76236 169910 76248
rect 170306 76236 170312 76248
rect 170364 76236 170370 76288
rect 171796 76276 171824 76384
rect 172698 76372 172704 76424
rect 172756 76412 172762 76424
rect 173342 76412 173348 76424
rect 172756 76384 173348 76412
rect 172756 76372 172762 76384
rect 173342 76372 173348 76384
rect 173400 76372 173406 76424
rect 172790 76304 172796 76356
rect 172848 76344 172854 76356
rect 173526 76344 173532 76356
rect 172848 76316 173532 76344
rect 172848 76304 172854 76316
rect 173526 76304 173532 76316
rect 173584 76304 173590 76356
rect 179138 76276 179144 76288
rect 171796 76248 179144 76276
rect 179138 76236 179144 76248
rect 179196 76236 179202 76288
rect 153286 76168 153292 76220
rect 153344 76208 153350 76220
rect 153838 76208 153844 76220
rect 153344 76180 153844 76208
rect 153344 76168 153350 76180
rect 153838 76168 153844 76180
rect 153896 76168 153902 76220
rect 168466 76168 168472 76220
rect 168524 76208 168530 76220
rect 175642 76208 175648 76220
rect 168524 76180 175648 76208
rect 168524 76168 168530 76180
rect 175642 76168 175648 76180
rect 175700 76168 175706 76220
rect 146386 76100 146392 76152
rect 146444 76140 146450 76152
rect 147214 76140 147220 76152
rect 146444 76112 147220 76140
rect 146444 76100 146450 76112
rect 147214 76100 147220 76112
rect 147272 76100 147278 76152
rect 157518 76100 157524 76152
rect 157576 76140 157582 76152
rect 179046 76140 179052 76152
rect 157576 76112 179052 76140
rect 157576 76100 157582 76112
rect 179046 76100 179052 76112
rect 179104 76100 179110 76152
rect 160370 76032 160376 76084
rect 160428 76072 160434 76084
rect 160554 76072 160560 76084
rect 160428 76044 160560 76072
rect 160428 76032 160434 76044
rect 160554 76032 160560 76044
rect 160612 76032 160618 76084
rect 168650 76032 168656 76084
rect 168708 76072 168714 76084
rect 170950 76072 170956 76084
rect 168708 76044 170956 76072
rect 168708 76032 168714 76044
rect 170950 76032 170956 76044
rect 171008 76032 171014 76084
rect 171502 76032 171508 76084
rect 171560 76072 171566 76084
rect 172146 76072 172152 76084
rect 171560 76044 172152 76072
rect 171560 76032 171566 76044
rect 172146 76032 172152 76044
rect 172204 76032 172210 76084
rect 141418 75964 141424 76016
rect 141476 76004 141482 76016
rect 141602 76004 141608 76016
rect 141476 75976 141608 76004
rect 141476 75964 141482 75976
rect 141602 75964 141608 75976
rect 141660 75964 141666 76016
rect 150618 75964 150624 76016
rect 150676 76004 150682 76016
rect 151354 76004 151360 76016
rect 150676 75976 151360 76004
rect 150676 75964 150682 75976
rect 151354 75964 151360 75976
rect 151412 75964 151418 76016
rect 151998 75964 152004 76016
rect 152056 76004 152062 76016
rect 152734 76004 152740 76016
rect 152056 75976 152740 76004
rect 152056 75964 152062 75976
rect 152734 75964 152740 75976
rect 152792 75964 152798 76016
rect 153010 75964 153016 76016
rect 153068 76004 153074 76016
rect 153930 76004 153936 76016
rect 153068 75976 153936 76004
rect 153068 75964 153074 75976
rect 153930 75964 153936 75976
rect 153988 75964 153994 76016
rect 166994 75964 167000 76016
rect 167052 76004 167058 76016
rect 176010 76004 176016 76016
rect 167052 75976 176016 76004
rect 167052 75964 167058 75976
rect 176010 75964 176016 75976
rect 176068 75964 176074 76016
rect 129090 75896 129096 75948
rect 129148 75936 129154 75948
rect 133598 75936 133604 75948
rect 129148 75908 133604 75936
rect 129148 75896 129154 75908
rect 133598 75896 133604 75908
rect 133656 75896 133662 75948
rect 138014 75896 138020 75948
rect 138072 75936 138078 75948
rect 141326 75936 141332 75948
rect 138072 75908 141332 75936
rect 138072 75896 138078 75908
rect 141326 75896 141332 75908
rect 141384 75896 141390 75948
rect 149054 75896 149060 75948
rect 149112 75936 149118 75948
rect 149238 75936 149244 75948
rect 149112 75908 149244 75936
rect 149112 75896 149118 75908
rect 149238 75896 149244 75908
rect 149296 75896 149302 75948
rect 150802 75896 150808 75948
rect 150860 75936 150866 75948
rect 151170 75936 151176 75948
rect 150860 75908 151176 75936
rect 150860 75896 150866 75908
rect 151170 75896 151176 75908
rect 151228 75896 151234 75948
rect 151722 75896 151728 75948
rect 151780 75936 151786 75948
rect 152458 75936 152464 75948
rect 151780 75908 152464 75936
rect 151780 75896 151786 75908
rect 152458 75896 152464 75908
rect 152516 75896 152522 75948
rect 153194 75896 153200 75948
rect 153252 75936 153258 75948
rect 154206 75936 154212 75948
rect 153252 75908 154212 75936
rect 153252 75896 153258 75908
rect 154206 75896 154212 75908
rect 154264 75896 154270 75948
rect 155034 75896 155040 75948
rect 155092 75936 155098 75948
rect 158530 75936 158536 75948
rect 155092 75908 158536 75936
rect 155092 75896 155098 75908
rect 158530 75896 158536 75908
rect 158588 75896 158594 75948
rect 159726 75896 159732 75948
rect 159784 75936 159790 75948
rect 159910 75936 159916 75948
rect 159784 75908 159916 75936
rect 159784 75896 159790 75908
rect 159910 75896 159916 75908
rect 159968 75896 159974 75948
rect 166534 75896 166540 75948
rect 166592 75936 166598 75948
rect 166718 75936 166724 75948
rect 166592 75908 166724 75936
rect 166592 75896 166598 75908
rect 166718 75896 166724 75908
rect 166776 75896 166782 75948
rect 168466 75896 168472 75948
rect 168524 75936 168530 75948
rect 168926 75936 168932 75948
rect 168524 75908 168932 75936
rect 168524 75896 168530 75908
rect 168926 75896 168932 75908
rect 168984 75896 168990 75948
rect 169110 75896 169116 75948
rect 169168 75936 169174 75948
rect 169662 75936 169668 75948
rect 169168 75908 169668 75936
rect 169168 75896 169174 75908
rect 169662 75896 169668 75908
rect 169720 75896 169726 75948
rect 170306 75896 170312 75948
rect 170364 75936 170370 75948
rect 170766 75936 170772 75948
rect 170364 75908 170772 75936
rect 170364 75896 170370 75908
rect 170766 75896 170772 75908
rect 170824 75896 170830 75948
rect 171134 75896 171140 75948
rect 171192 75936 171198 75948
rect 171686 75936 171692 75948
rect 171192 75908 171692 75936
rect 171192 75896 171198 75908
rect 171686 75896 171692 75908
rect 171744 75896 171750 75948
rect 118510 75828 118516 75880
rect 118568 75868 118574 75880
rect 580902 75868 580908 75880
rect 118568 75840 580908 75868
rect 118568 75828 118574 75840
rect 580902 75828 580908 75840
rect 580960 75828 580966 75880
rect 141326 75760 141332 75812
rect 141384 75800 141390 75812
rect 141786 75800 141792 75812
rect 141384 75772 141792 75800
rect 141384 75760 141390 75772
rect 141786 75760 141792 75772
rect 141844 75760 141850 75812
rect 145926 75760 145932 75812
rect 145984 75800 145990 75812
rect 191834 75800 191840 75812
rect 145984 75772 191840 75800
rect 145984 75760 145990 75772
rect 191834 75760 191840 75772
rect 191892 75760 191898 75812
rect 280338 75760 280344 75812
rect 280396 75800 280402 75812
rect 283190 75800 283196 75812
rect 280396 75772 283196 75800
rect 280396 75760 280402 75772
rect 283190 75760 283196 75772
rect 283248 75760 283254 75812
rect 148962 75692 148968 75744
rect 149020 75732 149026 75744
rect 220814 75732 220820 75744
rect 149020 75704 220820 75732
rect 149020 75692 149026 75704
rect 220814 75692 220820 75704
rect 220872 75692 220878 75744
rect 144638 75624 144644 75676
rect 144696 75664 144702 75676
rect 176194 75664 176200 75676
rect 144696 75636 176200 75664
rect 144696 75624 144702 75636
rect 176194 75624 176200 75636
rect 176252 75624 176258 75676
rect 177758 75624 177764 75676
rect 177816 75664 177822 75676
rect 256694 75664 256700 75676
rect 177816 75636 256700 75664
rect 177816 75624 177822 75636
rect 256694 75624 256700 75636
rect 256752 75624 256758 75676
rect 131298 75556 131304 75608
rect 131356 75596 131362 75608
rect 136174 75596 136180 75608
rect 131356 75568 136180 75596
rect 131356 75556 131362 75568
rect 136174 75556 136180 75568
rect 136232 75556 136238 75608
rect 153194 75556 153200 75608
rect 153252 75596 153258 75608
rect 154022 75596 154028 75608
rect 153252 75568 154028 75596
rect 153252 75556 153258 75568
rect 154022 75556 154028 75568
rect 154080 75556 154086 75608
rect 157702 75556 157708 75608
rect 157760 75596 157766 75608
rect 159726 75596 159732 75608
rect 157760 75568 159732 75596
rect 157760 75556 157766 75568
rect 159726 75556 159732 75568
rect 159784 75556 159790 75608
rect 159818 75556 159824 75608
rect 159876 75596 159882 75608
rect 262858 75596 262864 75608
rect 159876 75568 262864 75596
rect 159876 75556 159882 75568
rect 262858 75556 262864 75568
rect 262916 75556 262922 75608
rect 130930 75488 130936 75540
rect 130988 75528 130994 75540
rect 140590 75528 140596 75540
rect 130988 75500 140596 75528
rect 130988 75488 130994 75500
rect 140590 75488 140596 75500
rect 140648 75488 140654 75540
rect 151906 75488 151912 75540
rect 151964 75528 151970 75540
rect 274634 75528 274640 75540
rect 151964 75500 274640 75528
rect 151964 75488 151970 75500
rect 274634 75488 274640 75500
rect 274692 75488 274698 75540
rect 311894 75488 311900 75540
rect 311952 75528 311958 75540
rect 320542 75528 320548 75540
rect 311952 75500 320548 75528
rect 311952 75488 311958 75500
rect 320542 75488 320548 75500
rect 320600 75488 320606 75540
rect 127066 75420 127072 75472
rect 127124 75460 127130 75472
rect 140314 75460 140320 75472
rect 127124 75432 140320 75460
rect 127124 75420 127130 75432
rect 140314 75420 140320 75432
rect 140372 75420 140378 75472
rect 169202 75420 169208 75472
rect 169260 75460 169266 75472
rect 169260 75432 173664 75460
rect 169260 75420 169266 75432
rect 114554 75352 114560 75404
rect 114612 75392 114618 75404
rect 139118 75392 139124 75404
rect 114612 75364 139124 75392
rect 114612 75352 114618 75364
rect 139118 75352 139124 75364
rect 139176 75352 139182 75404
rect 159174 75352 159180 75404
rect 159232 75392 159238 75404
rect 159232 75364 165292 75392
rect 159232 75352 159238 75364
rect 137278 75284 137284 75336
rect 137336 75324 137342 75336
rect 157702 75324 157708 75336
rect 137336 75296 157708 75324
rect 137336 75284 137342 75296
rect 157702 75284 157708 75296
rect 157760 75284 157766 75336
rect 164326 75284 164332 75336
rect 164384 75324 164390 75336
rect 165062 75324 165068 75336
rect 164384 75296 165068 75324
rect 164384 75284 164390 75296
rect 165062 75284 165068 75296
rect 165120 75284 165126 75336
rect 75914 75216 75920 75268
rect 75972 75256 75978 75268
rect 131298 75256 131304 75268
rect 75972 75228 131304 75256
rect 75972 75216 75978 75228
rect 131298 75216 131304 75228
rect 131356 75216 131362 75268
rect 134242 75216 134248 75268
rect 134300 75256 134306 75268
rect 134702 75256 134708 75268
rect 134300 75228 134708 75256
rect 134300 75216 134306 75228
rect 134702 75216 134708 75228
rect 134760 75216 134766 75268
rect 135622 75216 135628 75268
rect 135680 75256 135686 75268
rect 136266 75256 136272 75268
rect 135680 75228 136272 75256
rect 135680 75216 135686 75228
rect 136266 75216 136272 75228
rect 136324 75216 136330 75268
rect 138382 75216 138388 75268
rect 138440 75256 138446 75268
rect 139302 75256 139308 75268
rect 138440 75228 139308 75256
rect 138440 75216 138446 75228
rect 139302 75216 139308 75228
rect 139360 75216 139366 75268
rect 139578 75216 139584 75268
rect 139636 75256 139642 75268
rect 140222 75256 140228 75268
rect 139636 75228 140228 75256
rect 139636 75216 139642 75228
rect 140222 75216 140228 75228
rect 140280 75216 140286 75268
rect 155310 75216 155316 75268
rect 155368 75256 155374 75268
rect 156874 75256 156880 75268
rect 155368 75228 156880 75256
rect 155368 75216 155374 75228
rect 156874 75216 156880 75228
rect 156932 75216 156938 75268
rect 161658 75216 161664 75268
rect 161716 75256 161722 75268
rect 161842 75256 161848 75268
rect 161716 75228 161848 75256
rect 161716 75216 161722 75228
rect 161842 75216 161848 75228
rect 161900 75216 161906 75268
rect 163130 75216 163136 75268
rect 163188 75256 163194 75268
rect 163498 75256 163504 75268
rect 163188 75228 163504 75256
rect 163188 75216 163194 75228
rect 163498 75216 163504 75228
rect 163556 75216 163562 75268
rect 164510 75216 164516 75268
rect 164568 75256 164574 75268
rect 164878 75256 164884 75268
rect 164568 75228 164884 75256
rect 164568 75216 164574 75228
rect 164878 75216 164884 75228
rect 164936 75216 164942 75268
rect 53834 75148 53840 75200
rect 53892 75188 53898 75200
rect 53892 75160 118694 75188
rect 53892 75148 53898 75160
rect 118666 75052 118694 75160
rect 134334 75148 134340 75200
rect 134392 75188 134398 75200
rect 135070 75188 135076 75200
rect 134392 75160 135076 75188
rect 134392 75148 134398 75160
rect 135070 75148 135076 75160
rect 135128 75148 135134 75200
rect 135714 75148 135720 75200
rect 135772 75188 135778 75200
rect 136542 75188 136548 75200
rect 135772 75160 136548 75188
rect 135772 75148 135778 75160
rect 136542 75148 136548 75160
rect 136600 75148 136606 75200
rect 162854 75148 162860 75200
rect 162912 75188 162918 75200
rect 163222 75188 163228 75200
rect 162912 75160 163228 75188
rect 162912 75148 162918 75160
rect 163222 75148 163228 75160
rect 163280 75148 163286 75200
rect 164602 75148 164608 75200
rect 164660 75188 164666 75200
rect 164970 75188 164976 75200
rect 164660 75160 164976 75188
rect 164660 75148 164666 75160
rect 164970 75148 164976 75160
rect 165028 75148 165034 75200
rect 131298 75080 131304 75132
rect 131356 75120 131362 75132
rect 132494 75120 132500 75132
rect 131356 75092 132500 75120
rect 131356 75080 131362 75092
rect 132494 75080 132500 75092
rect 132552 75080 132558 75132
rect 163130 75080 163136 75132
rect 163188 75120 163194 75132
rect 163774 75120 163780 75132
rect 163188 75092 163780 75120
rect 163188 75080 163194 75092
rect 163774 75080 163780 75092
rect 163832 75080 163838 75132
rect 164234 75080 164240 75132
rect 164292 75120 164298 75132
rect 165154 75120 165160 75132
rect 164292 75092 165160 75120
rect 164292 75080 164298 75092
rect 165154 75080 165160 75092
rect 165212 75080 165218 75132
rect 165264 75120 165292 75364
rect 166166 75352 166172 75404
rect 166224 75392 166230 75404
rect 166534 75392 166540 75404
rect 166224 75364 166540 75392
rect 166224 75352 166230 75364
rect 166534 75352 166540 75364
rect 166592 75352 166598 75404
rect 171134 75352 171140 75404
rect 171192 75392 171198 75404
rect 172054 75392 172060 75404
rect 171192 75364 172060 75392
rect 171192 75352 171198 75364
rect 172054 75352 172060 75364
rect 172112 75352 172118 75404
rect 173636 75392 173664 75432
rect 173802 75420 173808 75472
rect 173860 75460 173866 75472
rect 485774 75460 485780 75472
rect 173860 75432 485780 75460
rect 173860 75420 173866 75432
rect 485774 75420 485780 75432
rect 485832 75420 485838 75472
rect 496814 75392 496820 75404
rect 173636 75364 496820 75392
rect 496814 75352 496820 75364
rect 496872 75352 496878 75404
rect 165890 75284 165896 75336
rect 165948 75324 165954 75336
rect 166442 75324 166448 75336
rect 165948 75296 166448 75324
rect 165948 75284 165954 75296
rect 166442 75284 166448 75296
rect 166500 75284 166506 75336
rect 169386 75284 169392 75336
rect 169444 75324 169450 75336
rect 499574 75324 499580 75336
rect 169444 75296 499580 75324
rect 169444 75284 169450 75296
rect 499574 75284 499580 75296
rect 499632 75284 499638 75336
rect 165614 75216 165620 75268
rect 165672 75256 165678 75268
rect 166166 75256 166172 75268
rect 165672 75228 166172 75256
rect 165672 75216 165678 75228
rect 166166 75216 166172 75228
rect 166224 75216 166230 75268
rect 166994 75216 167000 75268
rect 167052 75256 167058 75268
rect 167822 75256 167828 75268
rect 167052 75228 167828 75256
rect 167052 75216 167058 75228
rect 167822 75216 167828 75228
rect 167880 75216 167886 75268
rect 170582 75216 170588 75268
rect 170640 75256 170646 75268
rect 514754 75256 514760 75268
rect 170640 75228 514760 75256
rect 170640 75216 170646 75228
rect 514754 75216 514760 75228
rect 514812 75216 514818 75268
rect 165798 75148 165804 75200
rect 165856 75188 165862 75200
rect 166258 75188 166264 75200
rect 165856 75160 166264 75188
rect 165856 75148 165862 75160
rect 166258 75148 166264 75160
rect 166316 75148 166322 75200
rect 175090 75188 175096 75200
rect 173452 75160 175096 75188
rect 173452 75120 173480 75160
rect 175090 75148 175096 75160
rect 175148 75148 175154 75200
rect 175918 75148 175924 75200
rect 175976 75188 175982 75200
rect 543734 75188 543740 75200
rect 175976 75160 543740 75188
rect 175976 75148 175982 75160
rect 543734 75148 543740 75160
rect 543792 75148 543798 75200
rect 165264 75092 173480 75120
rect 173894 75080 173900 75132
rect 173952 75120 173958 75132
rect 174446 75120 174452 75132
rect 173952 75092 174452 75120
rect 173952 75080 173958 75092
rect 174446 75080 174452 75092
rect 174504 75080 174510 75132
rect 134886 75052 134892 75064
rect 118666 75024 134892 75052
rect 134886 75012 134892 75024
rect 134944 75012 134950 75064
rect 160186 75012 160192 75064
rect 160244 75052 160250 75064
rect 160646 75052 160652 75064
rect 160244 75024 160652 75052
rect 160244 75012 160250 75024
rect 160646 75012 160652 75024
rect 160704 75012 160710 75064
rect 161566 75012 161572 75064
rect 161624 75052 161630 75064
rect 162118 75052 162124 75064
rect 161624 75024 162124 75052
rect 161624 75012 161630 75024
rect 162118 75012 162124 75024
rect 162176 75012 162182 75064
rect 163222 75012 163228 75064
rect 163280 75052 163286 75064
rect 163866 75052 163872 75064
rect 163280 75024 163872 75052
rect 163280 75012 163286 75024
rect 163866 75012 163872 75024
rect 163924 75012 163930 75064
rect 178126 75012 178132 75064
rect 178184 75052 178190 75064
rect 179230 75052 179236 75064
rect 178184 75024 179236 75052
rect 178184 75012 178190 75024
rect 179230 75012 179236 75024
rect 179288 75012 179294 75064
rect 142522 74944 142528 74996
rect 142580 74984 142586 74996
rect 142982 74984 142988 74996
rect 142580 74956 142988 74984
rect 142580 74944 142586 74956
rect 142982 74944 142988 74956
rect 143040 74944 143046 74996
rect 165154 74944 165160 74996
rect 165212 74984 165218 74996
rect 165430 74984 165436 74996
rect 165212 74956 165436 74984
rect 165212 74944 165218 74956
rect 165430 74944 165436 74956
rect 165488 74944 165494 74996
rect 160278 74740 160284 74792
rect 160336 74780 160342 74792
rect 160922 74780 160928 74792
rect 160336 74752 160928 74780
rect 160336 74740 160342 74752
rect 160922 74740 160928 74752
rect 160980 74740 160986 74792
rect 143810 74672 143816 74724
rect 143868 74712 143874 74724
rect 144178 74712 144184 74724
rect 143868 74684 144184 74712
rect 143868 74672 143874 74684
rect 144178 74672 144184 74684
rect 144236 74672 144242 74724
rect 168558 74672 168564 74724
rect 168616 74712 168622 74724
rect 169478 74712 169484 74724
rect 168616 74684 169484 74712
rect 168616 74672 168622 74684
rect 169478 74672 169484 74684
rect 169536 74672 169542 74724
rect 148594 74468 148600 74520
rect 148652 74508 148658 74520
rect 230474 74508 230480 74520
rect 148652 74480 230480 74508
rect 148652 74468 148658 74480
rect 230474 74468 230480 74480
rect 230532 74468 230538 74520
rect 157610 74400 157616 74452
rect 157668 74440 157674 74452
rect 242802 74440 242808 74452
rect 157668 74412 242808 74440
rect 157668 74400 157674 74412
rect 242802 74400 242808 74412
rect 242860 74400 242866 74452
rect 155494 74332 155500 74384
rect 155552 74372 155558 74384
rect 248966 74372 248972 74384
rect 155552 74344 248972 74372
rect 155552 74332 155558 74344
rect 248966 74332 248972 74344
rect 249024 74332 249030 74384
rect 93854 74264 93860 74316
rect 93912 74304 93918 74316
rect 137922 74304 137928 74316
rect 93912 74276 137928 74304
rect 93912 74264 93918 74276
rect 137922 74264 137928 74276
rect 137980 74264 137986 74316
rect 150158 74264 150164 74316
rect 150216 74304 150222 74316
rect 244366 74304 244372 74316
rect 150216 74276 244372 74304
rect 150216 74264 150222 74276
rect 244366 74264 244372 74276
rect 244424 74264 244430 74316
rect 89714 74196 89720 74248
rect 89772 74236 89778 74248
rect 137554 74236 137560 74248
rect 89772 74208 137560 74236
rect 89772 74196 89778 74208
rect 137554 74196 137560 74208
rect 137612 74196 137618 74248
rect 157610 74196 157616 74248
rect 157668 74236 157674 74248
rect 256786 74236 256792 74248
rect 157668 74208 256792 74236
rect 157668 74196 157674 74208
rect 256786 74196 256792 74208
rect 256844 74196 256850 74248
rect 86954 74128 86960 74180
rect 87012 74168 87018 74180
rect 137462 74168 137468 74180
rect 87012 74140 137468 74168
rect 87012 74128 87018 74140
rect 137462 74128 137468 74140
rect 137520 74128 137526 74180
rect 154666 74128 154672 74180
rect 154724 74168 154730 74180
rect 261478 74168 261484 74180
rect 154724 74140 261484 74168
rect 154724 74128 154730 74140
rect 261478 74128 261484 74140
rect 261536 74128 261542 74180
rect 57974 74060 57980 74112
rect 58032 74100 58038 74112
rect 134978 74100 134984 74112
rect 58032 74072 134984 74100
rect 58032 74060 58038 74072
rect 134978 74060 134984 74072
rect 135036 74060 135042 74112
rect 161106 74060 161112 74112
rect 161164 74100 161170 74112
rect 282178 74100 282184 74112
rect 161164 74072 282184 74100
rect 161164 74060 161170 74072
rect 282178 74060 282184 74072
rect 282236 74060 282242 74112
rect 51074 73992 51080 74044
rect 51132 74032 51138 74044
rect 134610 74032 134616 74044
rect 51132 74004 134616 74032
rect 51132 73992 51138 74004
rect 134610 73992 134616 74004
rect 134668 73992 134674 74044
rect 151906 73992 151912 74044
rect 151964 74032 151970 74044
rect 152550 74032 152556 74044
rect 151964 74004 152556 74032
rect 151964 73992 151970 74004
rect 152550 73992 152556 74004
rect 152608 73992 152614 74044
rect 157058 73992 157064 74044
rect 157116 74032 157122 74044
rect 281810 74032 281816 74044
rect 157116 74004 281816 74032
rect 157116 73992 157122 74004
rect 281810 73992 281816 74004
rect 281868 73992 281874 74044
rect 41414 73924 41420 73976
rect 41472 73964 41478 73976
rect 133782 73964 133788 73976
rect 41472 73936 133788 73964
rect 41472 73924 41478 73936
rect 133782 73924 133788 73936
rect 133840 73924 133846 73976
rect 158438 73924 158444 73976
rect 158496 73964 158502 73976
rect 290458 73964 290464 73976
rect 158496 73936 290464 73964
rect 158496 73924 158502 73936
rect 290458 73924 290464 73936
rect 290516 73924 290522 73976
rect 31754 73856 31760 73908
rect 31812 73896 31818 73908
rect 132126 73896 132132 73908
rect 31812 73868 132132 73896
rect 31812 73856 31818 73868
rect 132126 73856 132132 73868
rect 132184 73856 132190 73908
rect 155862 73856 155868 73908
rect 155920 73896 155926 73908
rect 295978 73896 295984 73908
rect 155920 73868 295984 73896
rect 155920 73856 155926 73868
rect 295978 73856 295984 73868
rect 296036 73856 296042 73908
rect 177298 73788 177304 73840
rect 177356 73828 177362 73840
rect 177666 73828 177672 73840
rect 177356 73800 177672 73828
rect 177356 73788 177362 73800
rect 177666 73788 177672 73800
rect 177724 73788 177730 73840
rect 178770 73788 178776 73840
rect 178828 73828 178834 73840
rect 446398 73828 446404 73840
rect 178828 73800 446404 73828
rect 178828 73788 178834 73800
rect 446398 73788 446404 73800
rect 446456 73788 446462 73840
rect 157610 73720 157616 73772
rect 157668 73760 157674 73772
rect 226518 73760 226524 73772
rect 157668 73732 226524 73760
rect 157668 73720 157674 73732
rect 226518 73720 226524 73732
rect 226576 73720 226582 73772
rect 132770 73652 132776 73704
rect 132828 73692 132834 73704
rect 133414 73692 133420 73704
rect 132828 73664 133420 73692
rect 132828 73652 132834 73664
rect 133414 73652 133420 73664
rect 133472 73652 133478 73704
rect 156230 73652 156236 73704
rect 156288 73692 156294 73704
rect 226426 73692 226432 73704
rect 156288 73664 226432 73692
rect 156288 73652 156294 73664
rect 226426 73652 226432 73664
rect 226484 73652 226490 73704
rect 158162 73584 158168 73636
rect 158220 73624 158226 73636
rect 178034 73624 178040 73636
rect 158220 73596 178040 73624
rect 158220 73584 158226 73596
rect 178034 73584 178040 73596
rect 178092 73584 178098 73636
rect 169018 73516 169024 73568
rect 169076 73556 169082 73568
rect 177298 73556 177304 73568
rect 169076 73528 177304 73556
rect 169076 73516 169082 73528
rect 177298 73516 177304 73528
rect 177356 73516 177362 73568
rect 170490 73448 170496 73500
rect 170548 73488 170554 73500
rect 177758 73488 177764 73500
rect 170548 73460 177764 73488
rect 170548 73448 170554 73460
rect 177758 73448 177764 73460
rect 177816 73448 177822 73500
rect 127618 73176 127624 73228
rect 127676 73216 127682 73228
rect 130286 73216 130292 73228
rect 127676 73188 130292 73216
rect 127676 73176 127682 73188
rect 130286 73176 130292 73188
rect 130344 73176 130350 73228
rect 136818 73176 136824 73228
rect 136876 73216 136882 73228
rect 141510 73216 141516 73228
rect 136876 73188 141516 73216
rect 136876 73176 136882 73188
rect 141510 73176 141516 73188
rect 141568 73176 141574 73228
rect 176102 73108 176108 73160
rect 176160 73148 176166 73160
rect 580166 73148 580172 73160
rect 176160 73120 580172 73148
rect 176160 73108 176166 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 156322 73040 156328 73092
rect 156380 73080 156386 73092
rect 255314 73080 255320 73092
rect 156380 73052 255320 73080
rect 156380 73040 156386 73052
rect 255314 73040 255320 73052
rect 255372 73040 255378 73092
rect 135990 73012 135996 73024
rect 118666 72984 135996 73012
rect 71774 72632 71780 72684
rect 71832 72672 71838 72684
rect 118666 72672 118694 72984
rect 135990 72972 135996 72984
rect 136048 72972 136054 73024
rect 175090 72972 175096 73024
rect 175148 73012 175154 73024
rect 281350 73012 281356 73024
rect 175148 72984 281356 73012
rect 175148 72972 175154 72984
rect 281350 72972 281356 72984
rect 281408 72972 281414 73024
rect 130930 72904 130936 72956
rect 130988 72904 130994 72956
rect 159726 72904 159732 72956
rect 159784 72944 159790 72956
rect 281442 72944 281448 72956
rect 159784 72916 281448 72944
rect 159784 72904 159790 72916
rect 281442 72904 281448 72916
rect 281500 72904 281506 72956
rect 130194 72700 130200 72752
rect 130252 72740 130258 72752
rect 130948 72740 130976 72904
rect 159542 72836 159548 72888
rect 159600 72876 159606 72888
rect 281994 72876 282000 72888
rect 159600 72848 282000 72876
rect 159600 72836 159606 72848
rect 281994 72836 282000 72848
rect 282052 72836 282058 72888
rect 159450 72768 159456 72820
rect 159508 72808 159514 72820
rect 281902 72808 281908 72820
rect 159508 72780 281908 72808
rect 159508 72768 159514 72780
rect 281902 72768 281908 72780
rect 281960 72768 281966 72820
rect 295334 72768 295340 72820
rect 295392 72808 295398 72820
rect 300302 72808 300308 72820
rect 295392 72780 300308 72808
rect 295392 72768 295398 72780
rect 300302 72768 300308 72780
rect 300360 72768 300366 72820
rect 130252 72712 130976 72740
rect 130252 72700 130258 72712
rect 158990 72700 158996 72752
rect 159048 72740 159054 72752
rect 299382 72740 299388 72752
rect 159048 72712 299388 72740
rect 159048 72700 159054 72712
rect 299382 72700 299388 72712
rect 299440 72700 299446 72752
rect 71832 72644 118694 72672
rect 71832 72632 71838 72644
rect 129826 72632 129832 72684
rect 129884 72672 129890 72684
rect 130470 72672 130476 72684
rect 129884 72644 130476 72672
rect 129884 72632 129890 72644
rect 130470 72632 130476 72644
rect 130528 72632 130534 72684
rect 158346 72632 158352 72684
rect 158404 72672 158410 72684
rect 311158 72672 311164 72684
rect 158404 72644 311164 72672
rect 158404 72632 158410 72644
rect 311158 72632 311164 72644
rect 311216 72632 311222 72684
rect 102134 72564 102140 72616
rect 102192 72604 102198 72616
rect 138934 72604 138940 72616
rect 102192 72576 138940 72604
rect 102192 72564 102198 72576
rect 138934 72564 138940 72576
rect 138992 72564 138998 72616
rect 165246 72564 165252 72616
rect 165304 72604 165310 72616
rect 347774 72604 347780 72616
rect 165304 72576 347780 72604
rect 165304 72564 165310 72576
rect 347774 72564 347780 72576
rect 347832 72564 347838 72616
rect 82814 72496 82820 72548
rect 82872 72536 82878 72548
rect 137738 72536 137744 72548
rect 82872 72508 137744 72536
rect 82872 72496 82878 72508
rect 137738 72496 137744 72508
rect 137796 72496 137802 72548
rect 159266 72496 159272 72548
rect 159324 72536 159330 72548
rect 349062 72536 349068 72548
rect 159324 72508 349068 72536
rect 159324 72496 159330 72508
rect 349062 72496 349068 72508
rect 349120 72496 349126 72548
rect 143166 72428 143172 72480
rect 143224 72468 143230 72480
rect 155954 72468 155960 72480
rect 143224 72440 155960 72468
rect 143224 72428 143230 72440
rect 155954 72428 155960 72440
rect 156012 72428 156018 72480
rect 167270 72428 167276 72480
rect 167328 72468 167334 72480
rect 417418 72468 417424 72480
rect 167328 72440 417424 72468
rect 167328 72428 167334 72440
rect 417418 72428 417424 72440
rect 417476 72428 417482 72480
rect 168374 72360 168380 72412
rect 168432 72400 168438 72412
rect 264974 72400 264980 72412
rect 168432 72372 264980 72400
rect 168432 72360 168438 72372
rect 264974 72360 264980 72372
rect 265032 72360 265038 72412
rect 178494 72292 178500 72344
rect 178552 72332 178558 72344
rect 275278 72332 275284 72344
rect 178552 72304 275284 72332
rect 178552 72292 178558 72304
rect 275278 72292 275284 72304
rect 275336 72292 275342 72344
rect 159082 72224 159088 72276
rect 159140 72264 159146 72276
rect 244274 72264 244280 72276
rect 159140 72236 244280 72264
rect 159140 72224 159146 72236
rect 244274 72224 244280 72236
rect 244332 72224 244338 72276
rect 135438 71748 135444 71800
rect 135496 71788 135502 71800
rect 141878 71788 141884 71800
rect 135496 71760 141884 71788
rect 135496 71748 135502 71760
rect 141878 71748 141884 71760
rect 141936 71748 141942 71800
rect 273530 71748 273536 71800
rect 273588 71788 273594 71800
rect 276014 71788 276020 71800
rect 273588 71760 276020 71788
rect 273588 71748 273594 71760
rect 276014 71748 276020 71760
rect 276072 71748 276078 71800
rect 283190 71680 283196 71732
rect 283248 71720 283254 71732
rect 289354 71720 289360 71732
rect 283248 71692 289360 71720
rect 283248 71680 283254 71692
rect 289354 71680 289360 71692
rect 289412 71680 289418 71732
rect 3418 71612 3424 71664
rect 3476 71652 3482 71664
rect 9030 71652 9036 71664
rect 3476 71624 9036 71652
rect 3476 71612 3482 71624
rect 9030 71612 9036 71624
rect 9088 71612 9094 71664
rect 179138 71612 179144 71664
rect 179196 71652 179202 71664
rect 195238 71652 195244 71664
rect 179196 71624 195244 71652
rect 179196 71612 179202 71624
rect 195238 71612 195244 71624
rect 195296 71612 195302 71664
rect 255314 71612 255320 71664
rect 255372 71652 255378 71664
rect 297358 71652 297364 71664
rect 255372 71624 297364 71652
rect 255372 71612 255378 71624
rect 297358 71612 297364 71624
rect 297416 71612 297422 71664
rect 154758 71544 154764 71596
rect 154816 71584 154822 71596
rect 257338 71584 257344 71596
rect 154816 71556 257344 71584
rect 154816 71544 154822 71556
rect 257338 71544 257344 71556
rect 257396 71544 257402 71596
rect 155218 71476 155224 71528
rect 155276 71516 155282 71528
rect 260190 71516 260196 71528
rect 155276 71488 260196 71516
rect 155276 71476 155282 71488
rect 260190 71476 260196 71488
rect 260248 71476 260254 71528
rect 155034 71408 155040 71460
rect 155092 71448 155098 71460
rect 272518 71448 272524 71460
rect 155092 71420 272524 71448
rect 155092 71408 155098 71420
rect 272518 71408 272524 71420
rect 272576 71408 272582 71460
rect 272886 71408 272892 71460
rect 272944 71448 272950 71460
rect 284294 71448 284300 71460
rect 272944 71420 284300 71448
rect 272944 71408 272950 71420
rect 284294 71408 284300 71420
rect 284352 71408 284358 71460
rect 156598 71340 156604 71392
rect 156656 71380 156662 71392
rect 280982 71380 280988 71392
rect 156656 71352 280988 71380
rect 156656 71340 156662 71352
rect 280982 71340 280988 71352
rect 281040 71340 281046 71392
rect 158898 71272 158904 71324
rect 158956 71312 158962 71324
rect 305730 71312 305736 71324
rect 158956 71284 305736 71312
rect 158956 71272 158962 71284
rect 305730 71272 305736 71284
rect 305788 71272 305794 71324
rect 318150 71272 318156 71324
rect 318208 71312 318214 71324
rect 332594 71312 332600 71324
rect 318208 71284 332600 71312
rect 318208 71272 318214 71284
rect 332594 71272 332600 71284
rect 332652 71272 332658 71324
rect 144730 71204 144736 71256
rect 144788 71244 144794 71256
rect 178310 71244 178316 71256
rect 144788 71216 178316 71244
rect 144788 71204 144794 71216
rect 178310 71204 178316 71216
rect 178368 71204 178374 71256
rect 179046 71204 179052 71256
rect 179104 71244 179110 71256
rect 334710 71244 334716 71256
rect 179104 71216 334716 71244
rect 179104 71204 179110 71216
rect 334710 71204 334716 71216
rect 334768 71204 334774 71256
rect 159910 71136 159916 71188
rect 159968 71176 159974 71188
rect 345658 71176 345664 71188
rect 159968 71148 345664 71176
rect 159968 71136 159974 71148
rect 345658 71136 345664 71148
rect 345716 71136 345722 71188
rect 167546 71068 167552 71120
rect 167604 71108 167610 71120
rect 456058 71108 456064 71120
rect 167604 71080 456064 71108
rect 167604 71068 167610 71080
rect 456058 71068 456064 71080
rect 456116 71068 456122 71120
rect 110414 71000 110420 71052
rect 110472 71040 110478 71052
rect 138566 71040 138572 71052
rect 110472 71012 138572 71040
rect 110472 71000 110478 71012
rect 138566 71000 138572 71012
rect 138624 71000 138630 71052
rect 167730 71000 167736 71052
rect 167788 71040 167794 71052
rect 467098 71040 467104 71052
rect 167788 71012 467104 71040
rect 167788 71000 167794 71012
rect 467098 71000 467104 71012
rect 467156 71000 467162 71052
rect 178034 70320 178040 70372
rect 178092 70360 178098 70372
rect 230842 70360 230848 70372
rect 178092 70332 230848 70360
rect 178092 70320 178098 70332
rect 230842 70320 230848 70332
rect 230900 70320 230906 70372
rect 156046 70252 156052 70304
rect 156104 70292 156110 70304
rect 226334 70292 226340 70304
rect 156104 70264 226340 70292
rect 156104 70252 156110 70264
rect 226334 70252 226340 70264
rect 226392 70252 226398 70304
rect 130838 70184 130844 70236
rect 130896 70224 130902 70236
rect 202322 70224 202328 70236
rect 130896 70196 202328 70224
rect 130896 70184 130902 70196
rect 202322 70184 202328 70196
rect 202380 70184 202386 70236
rect 226426 70184 226432 70236
rect 226484 70224 226490 70236
rect 273990 70224 273996 70236
rect 226484 70196 273996 70224
rect 226484 70184 226490 70196
rect 273990 70184 273996 70196
rect 274048 70184 274054 70236
rect 158530 70116 158536 70168
rect 158588 70156 158594 70168
rect 254578 70156 254584 70168
rect 158588 70128 254584 70156
rect 158588 70116 158594 70128
rect 254578 70116 254584 70128
rect 254636 70116 254642 70168
rect 256786 70116 256792 70168
rect 256844 70156 256850 70168
rect 280798 70156 280804 70168
rect 256844 70128 280804 70156
rect 256844 70116 256850 70128
rect 280798 70116 280804 70128
rect 280856 70116 280862 70168
rect 156966 70048 156972 70100
rect 157024 70088 157030 70100
rect 263042 70088 263048 70100
rect 157024 70060 263048 70088
rect 157024 70048 157030 70060
rect 263042 70048 263048 70060
rect 263100 70048 263106 70100
rect 310238 70048 310244 70100
rect 310296 70088 310302 70100
rect 312538 70088 312544 70100
rect 310296 70060 312544 70088
rect 310296 70048 310302 70060
rect 312538 70048 312544 70060
rect 312596 70048 312602 70100
rect 157702 69980 157708 70032
rect 157760 70020 157766 70032
rect 265618 70020 265624 70032
rect 157760 69992 265624 70020
rect 157760 69980 157766 69992
rect 265618 69980 265624 69992
rect 265676 69980 265682 70032
rect 155770 69912 155776 69964
rect 155828 69952 155834 69964
rect 271138 69952 271144 69964
rect 155828 69924 271144 69952
rect 155828 69912 155834 69924
rect 271138 69912 271144 69924
rect 271196 69912 271202 69964
rect 281350 69912 281356 69964
rect 281408 69952 281414 69964
rect 285766 69952 285772 69964
rect 281408 69924 285772 69952
rect 281408 69912 281414 69924
rect 285766 69912 285772 69924
rect 285824 69912 285830 69964
rect 299382 69912 299388 69964
rect 299440 69952 299446 69964
rect 309778 69952 309784 69964
rect 299440 69924 309784 69952
rect 299440 69912 299446 69924
rect 309778 69912 309784 69924
rect 309836 69912 309842 69964
rect 3418 69844 3424 69896
rect 3476 69884 3482 69896
rect 190730 69884 190736 69896
rect 3476 69856 190736 69884
rect 3476 69844 3482 69856
rect 190730 69844 190736 69856
rect 190788 69844 190794 69896
rect 244274 69844 244280 69896
rect 244332 69884 244338 69896
rect 349798 69884 349804 69896
rect 244332 69856 349804 69884
rect 244332 69844 244338 69856
rect 349798 69844 349804 69856
rect 349856 69844 349862 69896
rect 165338 69776 165344 69828
rect 165396 69816 165402 69828
rect 425054 69816 425060 69828
rect 165396 69788 425060 69816
rect 165396 69776 165402 69788
rect 425054 69776 425060 69788
rect 425112 69776 425118 69828
rect 446398 69776 446404 69828
rect 446456 69816 446462 69828
rect 460290 69816 460296 69828
rect 446456 69788 460296 69816
rect 446456 69776 446462 69788
rect 460290 69776 460296 69788
rect 460348 69776 460354 69828
rect 170398 69708 170404 69760
rect 170456 69748 170462 69760
rect 511994 69748 512000 69760
rect 170456 69720 512000 69748
rect 170456 69708 170462 69720
rect 511994 69708 512000 69720
rect 512052 69708 512058 69760
rect 2774 69640 2780 69692
rect 2832 69680 2838 69692
rect 130010 69680 130016 69692
rect 2832 69652 130016 69680
rect 2832 69640 2838 69652
rect 130010 69640 130016 69652
rect 130068 69640 130074 69692
rect 176470 69640 176476 69692
rect 176528 69680 176534 69692
rect 539594 69680 539600 69692
rect 176528 69652 539600 69680
rect 176528 69640 176534 69652
rect 539594 69640 539600 69652
rect 539652 69640 539658 69692
rect 178034 69572 178040 69624
rect 178092 69612 178098 69624
rect 178310 69612 178316 69624
rect 178092 69584 178316 69612
rect 178092 69572 178098 69584
rect 178310 69572 178316 69584
rect 178368 69572 178374 69624
rect 178862 69572 178868 69624
rect 178920 69612 178926 69624
rect 224954 69612 224960 69624
rect 178920 69584 224960 69612
rect 178920 69572 178926 69584
rect 224954 69572 224960 69584
rect 225012 69572 225018 69624
rect 226518 69572 226524 69624
rect 226576 69612 226582 69624
rect 274082 69612 274088 69624
rect 226576 69584 274088 69612
rect 226576 69572 226582 69584
rect 274082 69572 274088 69584
rect 274140 69572 274146 69624
rect 179414 69504 179420 69556
rect 179472 69544 179478 69556
rect 211062 69544 211068 69556
rect 179472 69516 211068 69544
rect 179472 69504 179478 69516
rect 211062 69504 211068 69516
rect 211120 69504 211126 69556
rect 310422 69504 310428 69556
rect 310480 69544 310486 69556
rect 318242 69544 318248 69556
rect 310480 69516 318248 69544
rect 310480 69504 310486 69516
rect 318242 69504 318248 69516
rect 318300 69504 318306 69556
rect 154666 69436 154672 69488
rect 154724 69476 154730 69488
rect 181990 69476 181996 69488
rect 154724 69448 181996 69476
rect 154724 69436 154730 69448
rect 181990 69436 181996 69448
rect 182048 69436 182054 69488
rect 281902 69232 281908 69284
rect 281960 69272 281966 69284
rect 284386 69272 284392 69284
rect 281960 69244 284392 69272
rect 281960 69232 281966 69244
rect 284386 69232 284392 69244
rect 284444 69232 284450 69284
rect 445478 69232 445484 69284
rect 445536 69272 445542 69284
rect 447134 69272 447140 69284
rect 445536 69244 447140 69272
rect 445536 69232 445542 69244
rect 447134 69232 447140 69244
rect 447192 69232 447198 69284
rect 281994 69164 282000 69216
rect 282052 69204 282058 69216
rect 284478 69204 284484 69216
rect 282052 69176 284484 69204
rect 282052 69164 282058 69176
rect 284478 69164 284484 69176
rect 284536 69164 284542 69216
rect 195238 68960 195244 69012
rect 195296 69000 195302 69012
rect 201126 69000 201132 69012
rect 195296 68972 201132 69000
rect 195296 68960 195302 68972
rect 201126 68960 201132 68972
rect 201184 68960 201190 69012
rect 281442 68960 281448 69012
rect 281500 69000 281506 69012
rect 298738 69000 298744 69012
rect 281500 68972 298744 69000
rect 281500 68960 281506 68972
rect 298738 68960 298744 68972
rect 298796 68960 298802 69012
rect 336734 68960 336740 69012
rect 336792 69000 336798 69012
rect 339494 69000 339500 69012
rect 336792 68972 339500 69000
rect 336792 68960 336798 68972
rect 339494 68960 339500 68972
rect 339552 68960 339558 69012
rect 222930 68892 222936 68944
rect 222988 68932 222994 68944
rect 294598 68932 294604 68944
rect 222988 68904 294604 68932
rect 222988 68892 222994 68904
rect 294598 68892 294604 68904
rect 294656 68892 294662 68944
rect 145558 68824 145564 68876
rect 145616 68864 145622 68876
rect 193214 68864 193220 68876
rect 145616 68836 193220 68864
rect 145616 68824 145622 68836
rect 193214 68824 193220 68836
rect 193272 68824 193278 68876
rect 242802 68824 242808 68876
rect 242860 68864 242866 68876
rect 318058 68864 318064 68876
rect 242860 68836 318064 68864
rect 242860 68824 242866 68836
rect 318058 68824 318064 68836
rect 318116 68824 318122 68876
rect 156874 68756 156880 68808
rect 156932 68796 156938 68808
rect 269850 68796 269856 68808
rect 156932 68768 269856 68796
rect 156932 68756 156938 68768
rect 269850 68756 269856 68768
rect 269908 68756 269914 68808
rect 281810 68756 281816 68808
rect 281868 68796 281874 68808
rect 316678 68796 316684 68808
rect 281868 68768 316684 68796
rect 281868 68756 281874 68768
rect 316678 68756 316684 68768
rect 316736 68756 316742 68808
rect 178954 68688 178960 68740
rect 179012 68728 179018 68740
rect 300394 68728 300400 68740
rect 179012 68700 300400 68728
rect 179012 68688 179018 68700
rect 300394 68688 300400 68700
rect 300452 68688 300458 68740
rect 332594 68688 332600 68740
rect 332652 68728 332658 68740
rect 340138 68728 340144 68740
rect 332652 68700 340144 68728
rect 332652 68688 332658 68700
rect 340138 68688 340144 68700
rect 340196 68688 340202 68740
rect 159634 68620 159640 68672
rect 159692 68660 159698 68672
rect 303154 68660 303160 68672
rect 159692 68632 303160 68660
rect 159692 68620 159698 68632
rect 303154 68620 303160 68632
rect 303212 68620 303218 68672
rect 320542 68620 320548 68672
rect 320600 68660 320606 68672
rect 359550 68660 359556 68672
rect 320600 68632 359556 68660
rect 320600 68620 320606 68632
rect 359550 68620 359556 68632
rect 359608 68620 359614 68672
rect 167086 68552 167092 68604
rect 167144 68592 167150 68604
rect 407114 68592 407120 68604
rect 167144 68564 407120 68592
rect 167144 68552 167150 68564
rect 407114 68552 407120 68564
rect 407172 68552 407178 68604
rect 167178 68484 167184 68536
rect 167236 68524 167242 68536
rect 420178 68524 420184 68536
rect 167236 68496 420184 68524
rect 167236 68484 167242 68496
rect 420178 68484 420184 68496
rect 420236 68484 420242 68536
rect 167270 68416 167276 68468
rect 167328 68456 167334 68468
rect 460198 68456 460204 68468
rect 167328 68428 460204 68456
rect 167328 68416 167334 68428
rect 460198 68416 460204 68428
rect 460256 68416 460262 68468
rect 169202 68348 169208 68400
rect 169260 68388 169266 68400
rect 498194 68388 498200 68400
rect 169260 68360 498200 68388
rect 169260 68348 169266 68360
rect 498194 68348 498200 68360
rect 498252 68348 498258 68400
rect 170306 68280 170312 68332
rect 170364 68320 170370 68332
rect 514846 68320 514852 68332
rect 170364 68292 514852 68320
rect 170364 68280 170370 68292
rect 514846 68280 514852 68292
rect 514904 68280 514910 68332
rect 289354 68212 289360 68264
rect 289412 68252 289418 68264
rect 300486 68252 300492 68264
rect 289412 68224 300492 68252
rect 289412 68212 289418 68224
rect 300486 68212 300492 68224
rect 300544 68212 300550 68264
rect 142798 67532 142804 67584
rect 142856 67572 142862 67584
rect 145558 67572 145564 67584
rect 142856 67544 145564 67572
rect 142856 67532 142862 67544
rect 145558 67532 145564 67544
rect 145616 67532 145622 67584
rect 262858 67532 262864 67584
rect 262916 67572 262922 67584
rect 266998 67572 267004 67584
rect 262916 67544 267004 67572
rect 262916 67532 262922 67544
rect 266998 67532 267004 67544
rect 267056 67532 267062 67584
rect 248966 67328 248972 67380
rect 249024 67368 249030 67380
rect 259546 67368 259552 67380
rect 249024 67340 259552 67368
rect 249024 67328 249030 67340
rect 259546 67328 259552 67340
rect 259604 67328 259610 67380
rect 264974 67328 264980 67380
rect 265032 67368 265038 67380
rect 273438 67368 273444 67380
rect 265032 67340 273444 67368
rect 265032 67328 265038 67340
rect 273438 67328 273444 67340
rect 273496 67328 273502 67380
rect 226334 67260 226340 67312
rect 226392 67300 226398 67312
rect 279418 67300 279424 67312
rect 226392 67272 279424 67300
rect 226392 67260 226398 67272
rect 279418 67260 279424 67272
rect 279476 67260 279482 67312
rect 211062 67192 211068 67244
rect 211120 67232 211126 67244
rect 269114 67232 269120 67244
rect 211120 67204 269120 67232
rect 211120 67192 211126 67204
rect 269114 67192 269120 67204
rect 269172 67192 269178 67244
rect 230842 67124 230848 67176
rect 230900 67164 230906 67176
rect 318150 67164 318156 67176
rect 230900 67136 318156 67164
rect 230900 67124 230906 67136
rect 318150 67124 318156 67136
rect 318208 67124 318214 67176
rect 181990 67056 181996 67108
rect 182048 67096 182054 67108
rect 285674 67096 285680 67108
rect 182048 67068 285680 67096
rect 182048 67056 182054 67068
rect 285674 67056 285680 67068
rect 285732 67056 285738 67108
rect 158254 66988 158260 67040
rect 158312 67028 158318 67040
rect 271598 67028 271604 67040
rect 158312 67000 271604 67028
rect 158312 66988 158318 67000
rect 271598 66988 271604 67000
rect 271656 66988 271662 67040
rect 276014 66988 276020 67040
rect 276072 67028 276078 67040
rect 282270 67028 282276 67040
rect 276072 67000 282276 67028
rect 276072 66988 276078 67000
rect 282270 66988 282276 67000
rect 282328 66988 282334 67040
rect 284294 66988 284300 67040
rect 284352 67028 284358 67040
rect 302970 67028 302976 67040
rect 284352 67000 302976 67028
rect 284352 66988 284358 67000
rect 302970 66988 302976 67000
rect 303028 66988 303034 67040
rect 224954 66920 224960 66972
rect 225012 66960 225018 66972
rect 348694 66960 348700 66972
rect 225012 66932 348700 66960
rect 225012 66920 225018 66932
rect 348694 66920 348700 66932
rect 348752 66920 348758 66972
rect 2866 66852 2872 66904
rect 2924 66892 2930 66904
rect 129918 66892 129924 66904
rect 2924 66864 129924 66892
rect 2924 66852 2930 66864
rect 129918 66852 129924 66864
rect 129976 66852 129982 66904
rect 164786 66852 164792 66904
rect 164844 66892 164850 66904
rect 437474 66892 437480 66904
rect 164844 66864 437480 66892
rect 164844 66852 164850 66864
rect 437474 66852 437480 66864
rect 437532 66852 437538 66904
rect 201126 66172 201132 66224
rect 201184 66212 201190 66224
rect 203518 66212 203524 66224
rect 201184 66184 203524 66212
rect 201184 66172 201190 66184
rect 203518 66172 203524 66184
rect 203576 66172 203582 66224
rect 260190 66172 260196 66224
rect 260248 66212 260254 66224
rect 263502 66212 263508 66224
rect 260248 66184 263508 66212
rect 260248 66172 260254 66184
rect 263502 66172 263508 66184
rect 263560 66172 263566 66224
rect 407114 66172 407120 66224
rect 407172 66212 407178 66224
rect 410518 66212 410524 66224
rect 407172 66184 410524 66212
rect 407172 66172 407178 66184
rect 410518 66172 410524 66184
rect 410576 66172 410582 66224
rect 447134 66172 447140 66224
rect 447192 66212 447198 66224
rect 450630 66212 450636 66224
rect 447192 66184 450636 66212
rect 447192 66172 447198 66184
rect 450630 66172 450636 66184
rect 450688 66172 450694 66224
rect 202322 66104 202328 66156
rect 202380 66144 202386 66156
rect 205358 66144 205364 66156
rect 202380 66116 205364 66144
rect 202380 66104 202386 66116
rect 205358 66104 205364 66116
rect 205416 66104 205422 66156
rect 339494 65764 339500 65816
rect 339552 65804 339558 65816
rect 345750 65804 345756 65816
rect 339552 65776 345756 65804
rect 339552 65764 339558 65776
rect 345750 65764 345756 65776
rect 345808 65764 345814 65816
rect 284386 65628 284392 65680
rect 284444 65668 284450 65680
rect 300118 65668 300124 65680
rect 284444 65640 300124 65668
rect 284444 65628 284450 65640
rect 300118 65628 300124 65640
rect 300176 65628 300182 65680
rect 284478 65560 284484 65612
rect 284536 65600 284542 65612
rect 300210 65600 300216 65612
rect 284536 65572 300216 65600
rect 284536 65560 284542 65572
rect 300210 65560 300216 65572
rect 300268 65560 300274 65612
rect 349062 65560 349068 65612
rect 349120 65600 349126 65612
rect 359458 65600 359464 65612
rect 349120 65572 359464 65600
rect 349120 65560 349126 65572
rect 359458 65560 359464 65572
rect 359516 65560 359522 65612
rect 164694 65492 164700 65544
rect 164752 65532 164758 65544
rect 434714 65532 434720 65544
rect 164752 65504 434720 65532
rect 164752 65492 164758 65504
rect 434714 65492 434720 65504
rect 434772 65492 434778 65544
rect 285766 64880 285772 64932
rect 285824 64920 285830 64932
rect 289078 64920 289084 64932
rect 285824 64892 289084 64920
rect 285824 64880 285830 64892
rect 289078 64880 289084 64892
rect 289136 64880 289142 64932
rect 294598 64336 294604 64388
rect 294656 64376 294662 64388
rect 301498 64376 301504 64388
rect 294656 64348 301504 64376
rect 294656 64336 294662 64348
rect 301498 64336 301504 64348
rect 301556 64336 301562 64388
rect 417418 64336 417424 64388
rect 417476 64376 417482 64388
rect 422938 64376 422944 64388
rect 417476 64348 422944 64376
rect 417476 64336 417482 64348
rect 422938 64336 422944 64348
rect 422996 64336 423002 64388
rect 285674 64268 285680 64320
rect 285732 64308 285738 64320
rect 294046 64308 294052 64320
rect 285732 64280 294052 64308
rect 285732 64268 285738 64280
rect 294046 64268 294052 64280
rect 294104 64268 294110 64320
rect 160646 64200 160652 64252
rect 160704 64240 160710 64252
rect 380894 64240 380900 64252
rect 160704 64212 380900 64240
rect 160704 64200 160710 64212
rect 380894 64200 380900 64212
rect 380952 64200 380958 64252
rect 174630 64132 174636 64184
rect 174688 64172 174694 64184
rect 568574 64172 568580 64184
rect 174688 64144 568580 64172
rect 174688 64132 174694 64144
rect 568574 64132 568580 64144
rect 568632 64132 568638 64184
rect 282270 64064 282276 64116
rect 282328 64104 282334 64116
rect 289354 64104 289360 64116
rect 282328 64076 289360 64104
rect 282328 64064 282334 64076
rect 289354 64064 289360 64076
rect 289412 64064 289418 64116
rect 254578 63996 254584 64048
rect 254636 64036 254642 64048
rect 260466 64036 260472 64048
rect 254636 64008 260472 64036
rect 254636 63996 254642 64008
rect 260466 63996 260472 64008
rect 260524 63996 260530 64048
rect 269114 63860 269120 63912
rect 269172 63900 269178 63912
rect 271874 63900 271880 63912
rect 269172 63872 271880 63900
rect 269172 63860 269178 63872
rect 271874 63860 271880 63872
rect 271932 63860 271938 63912
rect 263042 63724 263048 63776
rect 263100 63764 263106 63776
rect 265434 63764 265440 63776
rect 263100 63736 265440 63764
rect 263100 63724 263106 63736
rect 265434 63724 265440 63736
rect 265492 63724 265498 63776
rect 259546 63520 259552 63572
rect 259604 63560 259610 63572
rect 263410 63560 263416 63572
rect 259604 63532 263416 63560
rect 259604 63520 259610 63532
rect 263410 63520 263416 63532
rect 263468 63520 263474 63572
rect 282178 63452 282184 63504
rect 282236 63492 282242 63504
rect 287882 63492 287888 63504
rect 282236 63464 287888 63492
rect 282236 63452 282242 63464
rect 287882 63452 287888 63464
rect 287940 63452 287946 63504
rect 300394 63112 300400 63164
rect 300452 63152 300458 63164
rect 307662 63152 307668 63164
rect 300452 63124 307668 63152
rect 300452 63112 300458 63124
rect 307662 63112 307668 63124
rect 307720 63112 307726 63164
rect 300486 63044 300492 63096
rect 300544 63084 300550 63096
rect 303706 63084 303712 63096
rect 300544 63056 303712 63084
rect 300544 63044 300550 63056
rect 303706 63044 303712 63056
rect 303764 63044 303770 63096
rect 280982 62908 280988 62960
rect 281040 62948 281046 62960
rect 302326 62948 302332 62960
rect 281040 62920 302332 62948
rect 281040 62908 281046 62920
rect 302326 62908 302332 62920
rect 302384 62908 302390 62960
rect 261478 62840 261484 62892
rect 261536 62880 261542 62892
rect 276658 62880 276664 62892
rect 261536 62852 276664 62880
rect 261536 62840 261542 62852
rect 276658 62840 276664 62852
rect 276716 62840 276722 62892
rect 280890 62840 280896 62892
rect 280948 62880 280954 62892
rect 302234 62880 302240 62892
rect 280948 62852 302240 62880
rect 280948 62840 280954 62852
rect 302234 62840 302240 62852
rect 302292 62840 302298 62892
rect 460290 62840 460296 62892
rect 460348 62880 460354 62892
rect 464338 62880 464344 62892
rect 460348 62852 464344 62880
rect 460348 62840 460354 62852
rect 464338 62840 464344 62852
rect 464396 62840 464402 62892
rect 145466 62772 145472 62824
rect 145524 62812 145530 62824
rect 197354 62812 197360 62824
rect 145524 62784 197360 62812
rect 145524 62772 145530 62784
rect 197354 62772 197360 62784
rect 197412 62772 197418 62824
rect 261570 62772 261576 62824
rect 261628 62812 261634 62824
rect 284294 62812 284300 62824
rect 261628 62784 284300 62812
rect 261628 62772 261634 62784
rect 284294 62772 284300 62784
rect 284352 62772 284358 62824
rect 348694 62772 348700 62824
rect 348752 62812 348758 62824
rect 351914 62812 351920 62824
rect 348752 62784 351920 62812
rect 348752 62772 348758 62784
rect 351914 62772 351920 62784
rect 351972 62772 351978 62824
rect 439498 62772 439504 62824
rect 439556 62812 439562 62824
rect 463786 62812 463792 62824
rect 439556 62784 463792 62812
rect 439556 62772 439562 62784
rect 463786 62772 463792 62784
rect 463844 62772 463850 62824
rect 124214 62092 124220 62144
rect 124272 62132 124278 62144
rect 127710 62132 127716 62144
rect 124272 62104 127716 62132
rect 124272 62092 124278 62104
rect 127710 62092 127716 62104
rect 127768 62092 127774 62144
rect 297358 62092 297364 62144
rect 297416 62132 297422 62144
rect 302878 62132 302884 62144
rect 297416 62104 302884 62132
rect 297416 62092 297422 62104
rect 302878 62092 302884 62104
rect 302936 62092 302942 62144
rect 475378 62092 475384 62144
rect 475436 62132 475442 62144
rect 479518 62132 479524 62144
rect 475436 62104 479524 62132
rect 475436 62092 475442 62104
rect 479518 62092 479524 62104
rect 479576 62092 479582 62144
rect 271598 62024 271604 62076
rect 271656 62064 271662 62076
rect 277946 62064 277952 62076
rect 271656 62036 277952 62064
rect 271656 62024 271662 62036
rect 277946 62024 277952 62036
rect 278004 62024 278010 62076
rect 280798 62024 280804 62076
rect 280856 62064 280862 62076
rect 287698 62064 287704 62076
rect 280856 62036 287704 62064
rect 280856 62024 280862 62036
rect 287698 62024 287704 62036
rect 287756 62024 287762 62076
rect 311158 61888 311164 61940
rect 311216 61928 311222 61940
rect 315298 61928 315304 61940
rect 311216 61900 315304 61928
rect 311216 61888 311222 61900
rect 315298 61888 315304 61900
rect 315356 61888 315362 61940
rect 340138 61684 340144 61736
rect 340196 61724 340202 61736
rect 344278 61724 344284 61736
rect 340196 61696 344284 61724
rect 340196 61684 340202 61696
rect 344278 61684 344284 61696
rect 344336 61684 344342 61736
rect 359550 61412 359556 61464
rect 359608 61452 359614 61464
rect 361666 61452 361672 61464
rect 359608 61424 361672 61452
rect 359608 61412 359614 61424
rect 361666 61412 361672 61424
rect 361724 61412 361730 61464
rect 7558 61344 7564 61396
rect 7616 61384 7622 61396
rect 130102 61384 130108 61396
rect 7616 61356 130108 61384
rect 7616 61344 7622 61356
rect 130102 61344 130108 61356
rect 130160 61344 130166 61396
rect 301498 61344 301504 61396
rect 301556 61384 301562 61396
rect 313918 61384 313924 61396
rect 301556 61356 313924 61384
rect 301556 61344 301562 61356
rect 313918 61344 313924 61356
rect 313976 61344 313982 61396
rect 318242 61344 318248 61396
rect 318300 61384 318306 61396
rect 334618 61384 334624 61396
rect 318300 61356 334624 61384
rect 318300 61344 318306 61356
rect 334618 61344 334624 61356
rect 334676 61344 334682 61396
rect 289354 60800 289360 60852
rect 289412 60840 289418 60852
rect 291930 60840 291936 60852
rect 289412 60812 291936 60840
rect 289412 60800 289418 60812
rect 291930 60800 291936 60812
rect 291988 60800 291994 60852
rect 192570 60664 192576 60716
rect 192628 60704 192634 60716
rect 580166 60704 580172 60716
rect 192628 60676 580172 60704
rect 192628 60664 192634 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 265434 60596 265440 60648
rect 265492 60636 265498 60648
rect 269758 60636 269764 60648
rect 265492 60608 269764 60636
rect 265492 60596 265498 60608
rect 269758 60596 269764 60608
rect 269816 60596 269822 60648
rect 269850 60596 269856 60648
rect 269908 60636 269914 60648
rect 274726 60636 274732 60648
rect 269908 60608 274732 60636
rect 269908 60596 269914 60608
rect 274726 60596 274732 60608
rect 274784 60596 274790 60648
rect 142706 60460 142712 60512
rect 142764 60500 142770 60512
rect 148410 60500 148416 60512
rect 142764 60472 148416 60500
rect 142764 60460 142770 60472
rect 148410 60460 148416 60472
rect 148468 60460 148474 60512
rect 289170 60324 289176 60376
rect 289228 60364 289234 60376
rect 293954 60364 293960 60376
rect 289228 60336 293960 60364
rect 289228 60324 289234 60336
rect 293954 60324 293960 60336
rect 294012 60324 294018 60376
rect 312538 60256 312544 60308
rect 312596 60296 312602 60308
rect 315390 60296 315396 60308
rect 312596 60268 315396 60296
rect 312596 60256 312602 60268
rect 315390 60256 315396 60268
rect 315448 60256 315454 60308
rect 148318 60188 148324 60240
rect 148376 60228 148382 60240
rect 223574 60228 223580 60240
rect 148376 60200 223580 60228
rect 148376 60188 148382 60200
rect 223574 60188 223580 60200
rect 223632 60188 223638 60240
rect 257338 60188 257344 60240
rect 257396 60228 257402 60240
rect 261478 60228 261484 60240
rect 257396 60200 261484 60228
rect 257396 60188 257402 60200
rect 261478 60188 261484 60200
rect 261536 60188 261542 60240
rect 294046 60188 294052 60240
rect 294104 60228 294110 60240
rect 303062 60228 303068 60240
rect 294104 60200 303068 60228
rect 294104 60188 294110 60200
rect 303062 60188 303068 60200
rect 303120 60188 303126 60240
rect 303706 60188 303712 60240
rect 303764 60228 303770 60240
rect 326338 60228 326344 60240
rect 303764 60200 326344 60228
rect 303764 60188 303770 60200
rect 326338 60188 326344 60200
rect 326396 60188 326402 60240
rect 450630 60188 450636 60240
rect 450688 60228 450694 60240
rect 458818 60228 458824 60240
rect 450688 60200 458824 60228
rect 450688 60188 450694 60200
rect 458818 60188 458824 60200
rect 458876 60188 458882 60240
rect 168834 60120 168840 60172
rect 168892 60160 168898 60172
rect 491294 60160 491300 60172
rect 168892 60132 491300 60160
rect 168892 60120 168898 60132
rect 491294 60120 491300 60132
rect 491352 60120 491358 60172
rect 171870 60052 171876 60104
rect 171928 60092 171934 60104
rect 529934 60092 529940 60104
rect 171928 60064 529940 60092
rect 171928 60052 171934 60064
rect 529934 60052 529940 60064
rect 529992 60052 529998 60104
rect 117314 59984 117320 60036
rect 117372 60024 117378 60036
rect 129458 60024 129464 60036
rect 117372 59996 129464 60024
rect 117372 59984 117378 59996
rect 129458 59984 129464 59996
rect 129516 59984 129522 60036
rect 174538 59984 174544 60036
rect 174596 60024 174602 60036
rect 564434 60024 564440 60036
rect 174596 59996 564440 60024
rect 174596 59984 174602 59996
rect 564434 59984 564440 59996
rect 564492 59984 564498 60036
rect 302234 59712 302240 59764
rect 302292 59752 302298 59764
rect 306006 59752 306012 59764
rect 302292 59724 306012 59752
rect 302292 59712 302298 59724
rect 306006 59712 306012 59724
rect 306064 59712 306070 59764
rect 287882 59644 287888 59696
rect 287940 59684 287946 59696
rect 290550 59684 290556 59696
rect 287940 59656 290556 59684
rect 287940 59644 287946 59656
rect 290550 59644 290556 59656
rect 290608 59644 290614 59696
rect 302326 59576 302332 59628
rect 302384 59616 302390 59628
rect 306098 59616 306104 59628
rect 302384 59588 306104 59616
rect 302384 59576 302390 59588
rect 306098 59576 306104 59588
rect 306156 59576 306162 59628
rect 463786 59372 463792 59424
rect 463844 59412 463850 59424
rect 467190 59412 467196 59424
rect 463844 59384 467196 59412
rect 463844 59372 463850 59384
rect 467190 59372 467196 59384
rect 467248 59372 467254 59424
rect 205358 59304 205364 59356
rect 205416 59344 205422 59356
rect 210418 59344 210424 59356
rect 205416 59316 210424 59344
rect 205416 59304 205422 59316
rect 210418 59304 210424 59316
rect 210476 59304 210482 59356
rect 260466 59304 260472 59356
rect 260524 59344 260530 59356
rect 262214 59344 262220 59356
rect 260524 59316 262220 59344
rect 260524 59304 260530 59316
rect 262214 59304 262220 59316
rect 262272 59304 262278 59356
rect 263502 59304 263508 59356
rect 263560 59344 263566 59356
rect 268838 59344 268844 59356
rect 263560 59316 268844 59344
rect 263560 59304 263566 59316
rect 268838 59304 268844 59316
rect 268896 59304 268902 59356
rect 303246 59304 303252 59356
rect 303304 59344 303310 59356
rect 305822 59344 305828 59356
rect 303304 59316 305828 59344
rect 303304 59304 303310 59316
rect 305822 59304 305828 59316
rect 305880 59304 305886 59356
rect 334710 59304 334716 59356
rect 334768 59344 334774 59356
rect 337378 59344 337384 59356
rect 334768 59316 337384 59344
rect 334768 59304 334774 59316
rect 337378 59304 337384 59316
rect 337436 59304 337442 59356
rect 272518 58896 272524 58948
rect 272576 58936 272582 58948
rect 280982 58936 280988 58948
rect 272576 58908 280988 58936
rect 272576 58896 272582 58908
rect 280982 58896 280988 58908
rect 281040 58896 281046 58948
rect 271874 58828 271880 58880
rect 271932 58868 271938 58880
rect 286410 58868 286416 58880
rect 271932 58840 286416 58868
rect 271932 58828 271938 58840
rect 286410 58828 286416 58840
rect 286468 58828 286474 58880
rect 144178 58760 144184 58812
rect 144236 58800 144242 58812
rect 171870 58800 171876 58812
rect 144236 58772 171876 58800
rect 144236 58760 144242 58772
rect 171870 58760 171876 58772
rect 171928 58760 171934 58812
rect 273438 58760 273444 58812
rect 273496 58800 273502 58812
rect 283742 58800 283748 58812
rect 273496 58772 283748 58800
rect 273496 58760 273502 58772
rect 283742 58760 283748 58772
rect 283800 58760 283806 58812
rect 284294 58760 284300 58812
rect 284352 58800 284358 58812
rect 301314 58800 301320 58812
rect 284352 58772 301320 58800
rect 284352 58760 284358 58772
rect 301314 58760 301320 58772
rect 301372 58760 301378 58812
rect 351914 58760 351920 58812
rect 351972 58800 351978 58812
rect 369118 58800 369124 58812
rect 351972 58772 369124 58800
rect 351972 58760 351978 58772
rect 369118 58760 369124 58772
rect 369176 58760 369182 58812
rect 164602 58692 164608 58744
rect 164660 58732 164666 58744
rect 440234 58732 440240 58744
rect 164660 58704 440240 58732
rect 164660 58692 164666 58704
rect 440234 58692 440240 58704
rect 440292 58692 440298 58744
rect 102226 58624 102232 58676
rect 102284 58664 102290 58676
rect 130562 58664 130568 58676
rect 102284 58636 130568 58664
rect 102284 58624 102290 58636
rect 130562 58624 130568 58636
rect 130620 58624 130626 58676
rect 166994 58624 167000 58676
rect 167052 58664 167058 58676
rect 478874 58664 478880 58676
rect 167052 58636 478880 58664
rect 167052 58624 167058 58636
rect 478874 58624 478880 58636
rect 478932 58624 478938 58676
rect 277946 58556 277952 58608
rect 278004 58596 278010 58608
rect 283558 58596 283564 58608
rect 278004 58568 283564 58596
rect 278004 58556 278010 58568
rect 283558 58556 283564 58568
rect 283616 58556 283622 58608
rect 263410 57196 263416 57248
rect 263468 57236 263474 57248
rect 273254 57236 273260 57248
rect 263468 57208 273260 57236
rect 263468 57196 263474 57208
rect 273254 57196 273260 57208
rect 273312 57196 273318 57248
rect 279418 57196 279424 57248
rect 279476 57236 279482 57248
rect 287054 57236 287060 57248
rect 279476 57208 287060 57236
rect 279476 57196 279482 57208
rect 287054 57196 287060 57208
rect 287112 57196 287118 57248
rect 303154 57196 303160 57248
rect 303212 57236 303218 57248
rect 313182 57236 313188 57248
rect 303212 57208 313188 57236
rect 303212 57196 303218 57208
rect 313182 57196 313188 57208
rect 313240 57196 313246 57248
rect 460198 57196 460204 57248
rect 460256 57236 460262 57248
rect 464890 57236 464896 57248
rect 460256 57208 464896 57236
rect 460256 57196 460262 57208
rect 464890 57196 464896 57208
rect 464948 57196 464954 57248
rect 274726 56924 274732 56976
rect 274784 56964 274790 56976
rect 277762 56964 277768 56976
rect 274784 56936 277768 56964
rect 274784 56924 274790 56936
rect 277762 56924 277768 56936
rect 277820 56924 277826 56976
rect 262214 56516 262220 56568
rect 262272 56556 262278 56568
rect 266354 56556 266360 56568
rect 262272 56528 266360 56556
rect 262272 56516 262278 56528
rect 266354 56516 266360 56528
rect 266412 56516 266418 56568
rect 268838 56516 268844 56568
rect 268896 56556 268902 56568
rect 274266 56556 274272 56568
rect 268896 56528 274272 56556
rect 268896 56516 268902 56528
rect 274266 56516 274272 56528
rect 274324 56516 274330 56568
rect 280982 56516 280988 56568
rect 281040 56556 281046 56568
rect 286318 56556 286324 56568
rect 281040 56528 286324 56556
rect 281040 56516 281046 56528
rect 286318 56516 286324 56528
rect 286376 56516 286382 56568
rect 300302 56516 300308 56568
rect 300360 56556 300366 56568
rect 302234 56556 302240 56568
rect 300360 56528 302240 56556
rect 300360 56516 300366 56528
rect 302234 56516 302240 56528
rect 302292 56516 302298 56568
rect 309778 56516 309784 56568
rect 309836 56556 309842 56568
rect 314286 56556 314292 56568
rect 309836 56528 314292 56556
rect 309836 56516 309842 56528
rect 314286 56516 314292 56528
rect 314344 56516 314350 56568
rect 316678 56516 316684 56568
rect 316736 56556 316742 56568
rect 322198 56556 322204 56568
rect 316736 56528 322204 56556
rect 316736 56516 316742 56528
rect 322198 56516 322204 56528
rect 322256 56516 322262 56568
rect 301314 56448 301320 56500
rect 301372 56488 301378 56500
rect 305914 56488 305920 56500
rect 301372 56460 305920 56488
rect 301372 56448 301378 56460
rect 305914 56448 305920 56460
rect 305972 56448 305978 56500
rect 203518 55836 203524 55888
rect 203576 55876 203582 55888
rect 228358 55876 228364 55888
rect 203576 55848 228364 55876
rect 203576 55836 203582 55848
rect 228358 55836 228364 55848
rect 228416 55836 228422 55888
rect 271138 55836 271144 55888
rect 271196 55876 271202 55888
rect 291838 55876 291844 55888
rect 271196 55848 291844 55876
rect 271196 55836 271202 55848
rect 291838 55836 291844 55848
rect 291896 55836 291902 55888
rect 293954 55836 293960 55888
rect 294012 55876 294018 55888
rect 303522 55876 303528 55888
rect 294012 55848 303528 55876
rect 294012 55836 294018 55848
rect 303522 55836 303528 55848
rect 303580 55836 303586 55888
rect 307662 55836 307668 55888
rect 307720 55876 307726 55888
rect 321462 55876 321468 55888
rect 307720 55848 321468 55876
rect 307720 55836 307726 55848
rect 321462 55836 321468 55848
rect 321520 55836 321526 55888
rect 361666 55836 361672 55888
rect 361724 55876 361730 55888
rect 377398 55876 377404 55888
rect 361724 55848 377404 55876
rect 361724 55836 361730 55848
rect 377398 55836 377404 55848
rect 377456 55836 377462 55888
rect 306098 54748 306104 54800
rect 306156 54788 306162 54800
rect 309870 54788 309876 54800
rect 306156 54760 309876 54788
rect 306156 54748 306162 54760
rect 309870 54748 309876 54760
rect 309928 54748 309934 54800
rect 306006 54680 306012 54732
rect 306064 54720 306070 54732
rect 309778 54720 309784 54732
rect 306064 54692 309784 54720
rect 306064 54680 306070 54692
rect 309778 54680 309784 54692
rect 309836 54680 309842 54732
rect 305730 54612 305736 54664
rect 305788 54652 305794 54664
rect 312538 54652 312544 54664
rect 305788 54624 312544 54652
rect 305788 54612 305794 54624
rect 312538 54612 312544 54624
rect 312596 54612 312602 54664
rect 273254 54544 273260 54596
rect 273312 54584 273318 54596
rect 276106 54584 276112 54596
rect 273312 54556 276112 54584
rect 273312 54544 273318 54556
rect 276106 54544 276112 54556
rect 276164 54544 276170 54596
rect 305638 54544 305644 54596
rect 305696 54584 305702 54596
rect 323762 54584 323768 54596
rect 305696 54556 323768 54584
rect 305696 54544 305702 54556
rect 323762 54544 323768 54556
rect 323820 54544 323826 54596
rect 266998 54476 267004 54528
rect 267056 54516 267062 54528
rect 284294 54516 284300 54528
rect 267056 54488 284300 54516
rect 267056 54476 267062 54488
rect 284294 54476 284300 54488
rect 284352 54476 284358 54528
rect 287054 54476 287060 54528
rect 287112 54516 287118 54528
rect 319438 54516 319444 54528
rect 287112 54488 319444 54516
rect 287112 54476 287118 54488
rect 319438 54476 319444 54488
rect 319496 54476 319502 54528
rect 315390 54340 315396 54392
rect 315448 54380 315454 54392
rect 318334 54380 318340 54392
rect 315448 54352 318340 54380
rect 315448 54340 315454 54352
rect 318334 54340 318340 54352
rect 318392 54340 318398 54392
rect 291930 54136 291936 54188
rect 291988 54176 291994 54188
rect 299106 54176 299112 54188
rect 291988 54148 299112 54176
rect 291988 54136 291994 54148
rect 299106 54136 299112 54148
rect 299164 54136 299170 54188
rect 287698 54068 287704 54120
rect 287756 54108 287762 54120
rect 295334 54108 295340 54120
rect 287756 54080 295340 54108
rect 287756 54068 287762 54080
rect 295334 54068 295340 54080
rect 295392 54068 295398 54120
rect 410518 54068 410524 54120
rect 410576 54108 410582 54120
rect 413922 54108 413928 54120
rect 410576 54080 413928 54108
rect 410576 54068 410582 54080
rect 413922 54068 413928 54080
rect 413980 54068 413986 54120
rect 266354 53184 266360 53236
rect 266412 53224 266418 53236
rect 280798 53224 280804 53236
rect 266412 53196 280804 53224
rect 266412 53184 266418 53196
rect 280798 53184 280804 53196
rect 280856 53184 280862 53236
rect 295978 53184 295984 53236
rect 296036 53224 296042 53236
rect 309962 53224 309968 53236
rect 296036 53196 309968 53224
rect 296036 53184 296042 53196
rect 309962 53184 309968 53196
rect 310020 53184 310026 53236
rect 265618 53116 265624 53168
rect 265676 53156 265682 53168
rect 272518 53156 272524 53168
rect 265676 53128 272524 53156
rect 265676 53116 265682 53128
rect 272518 53116 272524 53128
rect 272576 53116 272582 53168
rect 274082 53116 274088 53168
rect 274140 53156 274146 53168
rect 297358 53156 297364 53168
rect 274140 53128 297364 53156
rect 274140 53116 274146 53128
rect 297358 53116 297364 53128
rect 297416 53116 297422 53168
rect 321462 53116 321468 53168
rect 321520 53156 321526 53168
rect 330478 53156 330484 53168
rect 321520 53128 330484 53156
rect 321520 53116 321526 53128
rect 330478 53116 330484 53128
rect 330536 53116 330542 53168
rect 261478 53048 261484 53100
rect 261536 53088 261542 53100
rect 273898 53088 273904 53100
rect 261536 53060 273904 53088
rect 261536 53048 261542 53060
rect 273898 53048 273904 53060
rect 273956 53048 273962 53100
rect 297450 53088 297456 53100
rect 277366 53060 297456 53088
rect 273990 52980 273996 53032
rect 274048 53020 274054 53032
rect 277366 53020 277394 53060
rect 297450 53048 297456 53060
rect 297508 53048 297514 53100
rect 326338 53048 326344 53100
rect 326396 53088 326402 53100
rect 350534 53088 350540 53100
rect 326396 53060 350540 53088
rect 326396 53048 326402 53060
rect 350534 53048 350540 53060
rect 350592 53048 350598 53100
rect 274048 52992 277394 53020
rect 274048 52980 274054 52992
rect 274266 52912 274272 52964
rect 274324 52952 274330 52964
rect 276014 52952 276020 52964
rect 274324 52924 276020 52952
rect 274324 52912 274330 52924
rect 276014 52912 276020 52924
rect 276072 52912 276078 52964
rect 302234 51960 302240 52012
rect 302292 52000 302298 52012
rect 304994 52000 305000 52012
rect 302292 51972 305000 52000
rect 302292 51960 302298 51972
rect 304994 51960 305000 51972
rect 305052 51960 305058 52012
rect 422938 51824 422944 51876
rect 422996 51864 423002 51876
rect 428458 51864 428464 51876
rect 422996 51836 428464 51864
rect 422996 51824 423002 51836
rect 428458 51824 428464 51836
rect 428516 51824 428522 51876
rect 315298 51756 315304 51808
rect 315356 51796 315362 51808
rect 320726 51796 320732 51808
rect 315356 51768 320732 51796
rect 315356 51756 315362 51768
rect 320726 51756 320732 51768
rect 320784 51756 320790 51808
rect 284294 51688 284300 51740
rect 284352 51728 284358 51740
rect 290826 51728 290832 51740
rect 284352 51700 290832 51728
rect 284352 51688 284358 51700
rect 290826 51688 290832 51700
rect 290884 51688 290890 51740
rect 303522 51688 303528 51740
rect 303580 51728 303586 51740
rect 311158 51728 311164 51740
rect 303580 51700 311164 51728
rect 303580 51688 303586 51700
rect 311158 51688 311164 51700
rect 311216 51688 311222 51740
rect 314286 51688 314292 51740
rect 314344 51728 314350 51740
rect 320818 51728 320824 51740
rect 314344 51700 320824 51728
rect 314344 51688 314350 51700
rect 320818 51688 320824 51700
rect 320876 51688 320882 51740
rect 210418 51620 210424 51672
rect 210476 51660 210482 51672
rect 212534 51660 212540 51672
rect 210476 51632 212540 51660
rect 210476 51620 210482 51632
rect 212534 51620 212540 51632
rect 212592 51620 212598 51672
rect 345750 51348 345756 51400
rect 345808 51388 345814 51400
rect 348418 51388 348424 51400
rect 345808 51360 348424 51388
rect 345808 51348 345814 51360
rect 348418 51348 348424 51360
rect 348476 51348 348482 51400
rect 330478 50804 330484 50856
rect 330536 50844 330542 50856
rect 336090 50844 336096 50856
rect 330536 50816 336096 50844
rect 330536 50804 330542 50816
rect 336090 50804 336096 50816
rect 336148 50804 336154 50856
rect 318150 50736 318156 50788
rect 318208 50776 318214 50788
rect 323670 50776 323676 50788
rect 318208 50748 323676 50776
rect 318208 50736 318214 50748
rect 323670 50736 323676 50748
rect 323728 50736 323734 50788
rect 290458 50532 290464 50584
rect 290516 50572 290522 50584
rect 293218 50572 293224 50584
rect 290516 50544 293224 50572
rect 290516 50532 290522 50544
rect 293218 50532 293224 50544
rect 293276 50532 293282 50584
rect 276014 50396 276020 50448
rect 276072 50436 276078 50448
rect 287606 50436 287612 50448
rect 276072 50408 287612 50436
rect 276072 50396 276078 50408
rect 287606 50396 287612 50408
rect 287664 50396 287670 50448
rect 305822 50396 305828 50448
rect 305880 50436 305886 50448
rect 310422 50436 310428 50448
rect 305880 50408 310428 50436
rect 305880 50396 305886 50408
rect 310422 50396 310428 50408
rect 310480 50396 310486 50448
rect 275278 50328 275284 50380
rect 275336 50368 275342 50380
rect 285674 50368 285680 50380
rect 275336 50340 285680 50368
rect 275336 50328 275342 50340
rect 285674 50328 285680 50340
rect 285732 50328 285738 50380
rect 290550 50328 290556 50380
rect 290608 50368 290614 50380
rect 305638 50368 305644 50380
rect 290608 50340 305644 50368
rect 290608 50328 290614 50340
rect 305638 50328 305644 50340
rect 305696 50328 305702 50380
rect 305914 50328 305920 50380
rect 305972 50368 305978 50380
rect 319530 50368 319536 50380
rect 305972 50340 319536 50368
rect 305972 50328 305978 50340
rect 319530 50328 319536 50340
rect 319588 50328 319594 50380
rect 299106 49784 299112 49836
rect 299164 49824 299170 49836
rect 301498 49824 301504 49836
rect 299164 49796 301504 49824
rect 299164 49784 299170 49796
rect 301498 49784 301504 49796
rect 301556 49784 301562 49836
rect 277762 49648 277768 49700
rect 277820 49688 277826 49700
rect 282914 49688 282920 49700
rect 277820 49660 282920 49688
rect 277820 49648 277826 49660
rect 282914 49648 282920 49660
rect 282972 49648 282978 49700
rect 313182 49648 313188 49700
rect 313240 49688 313246 49700
rect 318150 49688 318156 49700
rect 313240 49660 318156 49688
rect 313240 49648 313246 49660
rect 318150 49648 318156 49660
rect 318208 49648 318214 49700
rect 413922 49648 413928 49700
rect 413980 49688 413986 49700
rect 418154 49688 418160 49700
rect 413980 49660 418160 49688
rect 413980 49648 413986 49660
rect 418154 49648 418160 49660
rect 418212 49648 418218 49700
rect 464890 49648 464896 49700
rect 464948 49688 464954 49700
rect 471238 49688 471244 49700
rect 464948 49660 471244 49688
rect 464948 49648 464954 49660
rect 471238 49648 471244 49660
rect 471296 49648 471302 49700
rect 295334 49240 295340 49292
rect 295392 49280 295398 49292
rect 304258 49280 304264 49292
rect 295392 49252 304264 49280
rect 295392 49240 295398 49252
rect 304258 49240 304264 49252
rect 304316 49240 304322 49292
rect 300210 49172 300216 49224
rect 300268 49212 300274 49224
rect 310606 49212 310612 49224
rect 300268 49184 310612 49212
rect 300268 49172 300274 49184
rect 310606 49172 310612 49184
rect 310664 49172 310670 49224
rect 286410 49104 286416 49156
rect 286468 49144 286474 49156
rect 294598 49144 294604 49156
rect 286468 49116 294604 49144
rect 286468 49104 286474 49116
rect 294598 49104 294604 49116
rect 294656 49104 294662 49156
rect 300118 49104 300124 49156
rect 300176 49144 300182 49156
rect 310514 49144 310520 49156
rect 300176 49116 310520 49144
rect 300176 49104 300182 49116
rect 310514 49104 310520 49116
rect 310572 49104 310578 49156
rect 290826 49036 290832 49088
rect 290884 49076 290890 49088
rect 308490 49076 308496 49088
rect 290884 49048 308496 49076
rect 290884 49036 290890 49048
rect 308490 49036 308496 49048
rect 308548 49036 308554 49088
rect 177206 48968 177212 49020
rect 177264 49008 177270 49020
rect 440326 49008 440332 49020
rect 177264 48980 440332 49008
rect 177264 48968 177270 48980
rect 440326 48968 440332 48980
rect 440384 48968 440390 49020
rect 287606 48220 287612 48272
rect 287664 48260 287670 48272
rect 291930 48260 291936 48272
rect 287664 48232 291936 48260
rect 287664 48220 287670 48232
rect 291930 48220 291936 48232
rect 291988 48220 291994 48272
rect 318058 48220 318064 48272
rect 318116 48260 318122 48272
rect 323578 48260 323584 48272
rect 318116 48232 323584 48260
rect 318116 48220 318122 48232
rect 323578 48220 323584 48232
rect 323636 48220 323642 48272
rect 318334 48152 318340 48204
rect 318392 48192 318398 48204
rect 321002 48192 321008 48204
rect 318392 48164 321008 48192
rect 318392 48152 318398 48164
rect 321002 48152 321008 48164
rect 321060 48152 321066 48204
rect 276658 47676 276664 47728
rect 276716 47716 276722 47728
rect 282178 47716 282184 47728
rect 276716 47688 282184 47716
rect 276716 47676 276722 47688
rect 282178 47676 282184 47688
rect 282236 47676 282242 47728
rect 276106 47608 276112 47660
rect 276164 47648 276170 47660
rect 284938 47648 284944 47660
rect 276164 47620 284944 47648
rect 276164 47608 276170 47620
rect 284938 47608 284944 47620
rect 284996 47608 285002 47660
rect 269758 47540 269764 47592
rect 269816 47580 269822 47592
rect 283650 47580 283656 47592
rect 269816 47552 283656 47580
rect 269816 47540 269822 47552
rect 283650 47540 283656 47552
rect 283708 47540 283714 47592
rect 285674 47540 285680 47592
rect 285732 47580 285738 47592
rect 293862 47580 293868 47592
rect 285732 47552 293868 47580
rect 285732 47540 285738 47552
rect 293862 47540 293868 47552
rect 293920 47540 293926 47592
rect 304994 47540 305000 47592
rect 305052 47580 305058 47592
rect 309594 47580 309600 47592
rect 305052 47552 309600 47580
rect 305052 47540 305058 47552
rect 309594 47540 309600 47552
rect 309652 47540 309658 47592
rect 458818 47540 458824 47592
rect 458876 47580 458882 47592
rect 461302 47580 461308 47592
rect 458876 47552 461308 47580
rect 458876 47540 458882 47552
rect 461302 47540 461308 47552
rect 461360 47540 461366 47592
rect 467190 47540 467196 47592
rect 467248 47580 467254 47592
rect 476758 47580 476764 47592
rect 467248 47552 476764 47580
rect 467248 47540 467254 47552
rect 476758 47540 476764 47552
rect 476816 47540 476822 47592
rect 118418 46860 118424 46912
rect 118476 46900 118482 46912
rect 580166 46900 580172 46912
rect 118476 46872 580172 46900
rect 118476 46860 118482 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 310514 46792 310520 46844
rect 310572 46832 310578 46844
rect 313274 46832 313280 46844
rect 310572 46804 313280 46832
rect 310572 46792 310578 46804
rect 313274 46792 313280 46804
rect 313332 46792 313338 46844
rect 319438 46792 319444 46844
rect 319496 46832 319502 46844
rect 322842 46832 322848 46844
rect 319496 46804 322848 46832
rect 319496 46792 319502 46804
rect 322842 46792 322848 46804
rect 322900 46792 322906 46844
rect 310606 46724 310612 46776
rect 310664 46764 310670 46776
rect 313458 46764 313464 46776
rect 310664 46736 313464 46764
rect 310664 46724 310670 46736
rect 313458 46724 313464 46736
rect 313516 46724 313522 46776
rect 282914 46180 282920 46232
rect 282972 46220 282978 46232
rect 290642 46220 290648 46232
rect 282972 46192 290648 46220
rect 282972 46180 282978 46192
rect 290642 46180 290648 46192
rect 290700 46180 290706 46232
rect 303062 46180 303068 46232
rect 303120 46220 303126 46232
rect 308398 46220 308404 46232
rect 303120 46192 308404 46220
rect 303120 46180 303126 46192
rect 308398 46180 308404 46192
rect 308456 46180 308462 46232
rect 310422 46180 310428 46232
rect 310480 46220 310486 46232
rect 316770 46220 316776 46232
rect 310480 46192 316776 46220
rect 310480 46180 310486 46192
rect 316770 46180 316776 46192
rect 316828 46180 316834 46232
rect 320726 46180 320732 46232
rect 320784 46220 320790 46232
rect 338758 46220 338764 46232
rect 320784 46192 338764 46220
rect 320784 46180 320790 46192
rect 338758 46180 338764 46192
rect 338816 46180 338822 46232
rect 350534 46180 350540 46232
rect 350592 46220 350598 46232
rect 362218 46220 362224 46232
rect 350592 46192 362224 46220
rect 350592 46180 350598 46192
rect 362218 46180 362224 46192
rect 362276 46180 362282 46232
rect 418154 46180 418160 46232
rect 418212 46220 418218 46232
rect 429102 46220 429108 46232
rect 418212 46192 429108 46220
rect 418212 46180 418218 46192
rect 429102 46180 429108 46192
rect 429160 46180 429166 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 178218 45540 178224 45552
rect 3476 45512 178224 45540
rect 3476 45500 3482 45512
rect 178218 45500 178224 45512
rect 178276 45500 178282 45552
rect 284938 45500 284944 45552
rect 284996 45540 285002 45552
rect 287606 45540 287612 45552
rect 284996 45512 287612 45540
rect 284996 45500 285002 45512
rect 287606 45500 287612 45512
rect 287664 45500 287670 45552
rect 293862 44956 293868 45008
rect 293920 44996 293926 45008
rect 302234 44996 302240 45008
rect 293920 44968 302240 44996
rect 293920 44956 293926 44968
rect 302234 44956 302240 44968
rect 302292 44956 302298 45008
rect 228358 44888 228364 44940
rect 228416 44928 228422 44940
rect 233878 44928 233884 44940
rect 228416 44900 233884 44928
rect 228416 44888 228422 44900
rect 233878 44888 233884 44900
rect 233936 44888 233942 44940
rect 294598 44888 294604 44940
rect 294656 44928 294662 44940
rect 309042 44928 309048 44940
rect 294656 44900 309048 44928
rect 294656 44888 294662 44900
rect 309042 44888 309048 44900
rect 309100 44888 309106 44940
rect 175274 44820 175280 44872
rect 175332 44860 175338 44872
rect 580258 44860 580264 44872
rect 175332 44832 580264 44860
rect 175332 44820 175338 44832
rect 580258 44820 580264 44832
rect 580316 44820 580322 44872
rect 298738 44684 298744 44736
rect 298796 44724 298802 44736
rect 303798 44724 303804 44736
rect 298796 44696 303804 44724
rect 298796 44684 298802 44696
rect 303798 44684 303804 44696
rect 303856 44684 303862 44736
rect 311158 44548 311164 44600
rect 311216 44588 311222 44600
rect 317322 44588 317328 44600
rect 311216 44560 317328 44588
rect 311216 44548 311222 44560
rect 317322 44548 317328 44560
rect 317380 44548 317386 44600
rect 286318 44412 286324 44464
rect 286376 44452 286382 44464
rect 289722 44452 289728 44464
rect 286376 44424 289728 44452
rect 286376 44412 286382 44424
rect 289722 44412 289728 44424
rect 289780 44412 289786 44464
rect 320818 44276 320824 44328
rect 320876 44316 320882 44328
rect 323026 44316 323032 44328
rect 320876 44288 323032 44316
rect 320876 44276 320882 44288
rect 323026 44276 323032 44288
rect 323084 44276 323090 44328
rect 359458 43732 359464 43784
rect 359516 43772 359522 43784
rect 363598 43772 363604 43784
rect 359516 43744 363604 43772
rect 359516 43732 359522 43744
rect 363598 43732 363604 43744
rect 363656 43732 363662 43784
rect 308490 43528 308496 43580
rect 308548 43568 308554 43580
rect 317046 43568 317052 43580
rect 308548 43540 317052 43568
rect 308548 43528 308554 43540
rect 317046 43528 317052 43540
rect 317104 43528 317110 43580
rect 309962 43460 309968 43512
rect 310020 43500 310026 43512
rect 319438 43500 319444 43512
rect 310020 43472 319444 43500
rect 310020 43460 310026 43472
rect 319438 43460 319444 43472
rect 319496 43460 319502 43512
rect 323762 43460 323768 43512
rect 323820 43500 323826 43512
rect 326062 43500 326068 43512
rect 323820 43472 326068 43500
rect 323820 43460 323826 43472
rect 326062 43460 326068 43472
rect 326120 43460 326126 43512
rect 177942 43392 177948 43444
rect 178000 43432 178006 43444
rect 447134 43432 447140 43444
rect 178000 43404 447140 43432
rect 178000 43392 178006 43404
rect 447134 43392 447140 43404
rect 447192 43392 447198 43444
rect 309870 43324 309876 43376
rect 309928 43364 309934 43376
rect 312262 43364 312268 43376
rect 309928 43336 312268 43364
rect 309928 43324 309934 43336
rect 312262 43324 312268 43336
rect 312320 43324 312326 43376
rect 309778 43188 309784 43240
rect 309836 43228 309842 43240
rect 311894 43228 311900 43240
rect 309836 43200 311900 43228
rect 309836 43188 309842 43200
rect 311894 43188 311900 43200
rect 311952 43188 311958 43240
rect 456058 43052 456064 43104
rect 456116 43092 456122 43104
rect 458542 43092 458548 43104
rect 456116 43064 458548 43092
rect 456116 43052 456122 43064
rect 458542 43052 458548 43064
rect 458600 43052 458606 43104
rect 297450 42848 297456 42900
rect 297508 42888 297514 42900
rect 300762 42888 300768 42900
rect 297508 42860 300768 42888
rect 297508 42848 297514 42860
rect 300762 42848 300768 42860
rect 300820 42848 300826 42900
rect 297358 42780 297364 42832
rect 297416 42820 297422 42832
rect 300118 42820 300124 42832
rect 297416 42792 300124 42820
rect 297416 42780 297422 42792
rect 300118 42780 300124 42792
rect 300176 42780 300182 42832
rect 287606 42372 287612 42424
rect 287664 42412 287670 42424
rect 292022 42412 292028 42424
rect 287664 42384 292028 42412
rect 287664 42372 287670 42384
rect 292022 42372 292028 42384
rect 292080 42372 292086 42424
rect 289078 42100 289084 42152
rect 289136 42140 289142 42152
rect 297634 42140 297640 42152
rect 289136 42112 297640 42140
rect 289136 42100 289142 42112
rect 297634 42100 297640 42112
rect 297692 42100 297698 42152
rect 334618 42100 334624 42152
rect 334676 42140 334682 42152
rect 340138 42140 340144 42152
rect 334676 42112 340144 42140
rect 334676 42100 334682 42112
rect 340138 42100 340144 42112
rect 340196 42100 340202 42152
rect 293218 42032 293224 42084
rect 293276 42072 293282 42084
rect 303706 42072 303712 42084
rect 293276 42044 303712 42072
rect 293276 42032 293282 42044
rect 303706 42032 303712 42044
rect 303764 42032 303770 42084
rect 319530 42032 319536 42084
rect 319588 42072 319594 42084
rect 336182 42072 336188 42084
rect 319588 42044 336188 42072
rect 319588 42032 319594 42044
rect 336182 42032 336188 42044
rect 336240 42032 336246 42084
rect 322198 41556 322204 41608
rect 322256 41596 322262 41608
rect 324958 41596 324964 41608
rect 322256 41568 324964 41596
rect 322256 41556 322262 41568
rect 324958 41556 324964 41568
rect 325016 41556 325022 41608
rect 313918 41352 313924 41404
rect 313976 41392 313982 41404
rect 316678 41392 316684 41404
rect 313976 41364 316684 41392
rect 313976 41352 313982 41364
rect 316678 41352 316684 41364
rect 316736 41352 316742 41404
rect 322842 41352 322848 41404
rect 322900 41392 322906 41404
rect 327718 41392 327724 41404
rect 322900 41364 327724 41392
rect 322900 41352 322906 41364
rect 327718 41352 327724 41364
rect 327776 41352 327782 41404
rect 317322 41284 317328 41336
rect 317380 41324 317386 41336
rect 325050 41324 325056 41336
rect 317380 41296 325056 41324
rect 317380 41284 317386 41296
rect 325050 41284 325056 41296
rect 325108 41284 325114 41336
rect 309042 41216 309048 41268
rect 309100 41256 309106 41268
rect 310698 41256 310704 41268
rect 309100 41228 310704 41256
rect 309100 41216 309106 41228
rect 310698 41216 310704 41228
rect 310756 41216 310762 41268
rect 309594 40740 309600 40792
rect 309652 40780 309658 40792
rect 321094 40780 321100 40792
rect 309652 40752 321100 40780
rect 309652 40740 309658 40752
rect 321094 40740 321100 40752
rect 321152 40740 321158 40792
rect 99374 40672 99380 40724
rect 99432 40712 99438 40724
rect 130470 40712 130476 40724
rect 99432 40684 130476 40712
rect 99432 40672 99438 40684
rect 130470 40672 130476 40684
rect 130528 40672 130534 40724
rect 233878 40672 233884 40724
rect 233936 40712 233942 40724
rect 245654 40712 245660 40724
rect 233936 40684 245660 40712
rect 233936 40672 233942 40684
rect 245654 40672 245660 40684
rect 245712 40672 245718 40724
rect 305638 40672 305644 40724
rect 305696 40712 305702 40724
rect 322934 40712 322940 40724
rect 305696 40684 322940 40712
rect 305696 40672 305702 40684
rect 322934 40672 322940 40684
rect 322992 40672 322998 40724
rect 429102 40672 429108 40724
rect 429160 40712 429166 40724
rect 439498 40712 439504 40724
rect 429160 40684 439504 40712
rect 429160 40672 429166 40684
rect 439498 40672 439504 40684
rect 439556 40672 439562 40724
rect 290642 39992 290648 40044
rect 290700 40032 290706 40044
rect 294598 40032 294604 40044
rect 290700 40004 294604 40032
rect 290700 39992 290706 40004
rect 294598 39992 294604 40004
rect 294656 39992 294662 40044
rect 303706 39992 303712 40044
rect 303764 40032 303770 40044
rect 307018 40032 307024 40044
rect 303764 40004 307024 40032
rect 303764 39992 303770 40004
rect 307018 39992 307024 40004
rect 307076 39992 307082 40044
rect 313458 39992 313464 40044
rect 313516 40032 313522 40044
rect 317230 40032 317236 40044
rect 313516 40004 317236 40032
rect 313516 39992 313522 40004
rect 317230 39992 317236 40004
rect 317288 39992 317294 40044
rect 461302 39992 461308 40044
rect 461360 40032 461366 40044
rect 468478 40032 468484 40044
rect 461360 40004 468484 40032
rect 461360 39992 461366 40004
rect 468478 39992 468484 40004
rect 468536 39992 468542 40044
rect 313274 39924 313280 39976
rect 313332 39964 313338 39976
rect 317322 39964 317328 39976
rect 313332 39936 317328 39964
rect 313332 39924 313338 39936
rect 317322 39924 317328 39936
rect 317380 39924 317386 39976
rect 312262 39856 312268 39908
rect 312320 39896 312326 39908
rect 318518 39896 318524 39908
rect 312320 39868 318524 39896
rect 312320 39856 312326 39868
rect 318518 39856 318524 39868
rect 318576 39856 318582 39908
rect 311894 39788 311900 39840
rect 311952 39828 311958 39840
rect 318426 39828 318432 39840
rect 311952 39800 318432 39828
rect 311952 39788 311958 39800
rect 318426 39788 318432 39800
rect 318484 39788 318490 39840
rect 301498 39380 301504 39432
rect 301556 39420 301562 39432
rect 315298 39420 315304 39432
rect 301556 39392 315304 39420
rect 301556 39380 301562 39392
rect 315298 39380 315304 39392
rect 315356 39380 315362 39432
rect 318150 39380 318156 39432
rect 318208 39420 318214 39432
rect 337930 39420 337936 39432
rect 318208 39392 337936 39420
rect 318208 39380 318214 39392
rect 337930 39380 337936 39392
rect 337988 39380 337994 39432
rect 177850 39312 177856 39364
rect 177908 39352 177914 39364
rect 431954 39352 431960 39364
rect 177908 39324 431960 39352
rect 177908 39312 177914 39324
rect 431954 39312 431960 39324
rect 432012 39312 432018 39364
rect 338758 38428 338764 38480
rect 338816 38468 338822 38480
rect 347130 38468 347136 38480
rect 338816 38440 347136 38468
rect 338816 38428 338822 38440
rect 347130 38428 347136 38440
rect 347188 38428 347194 38480
rect 303798 37884 303804 37936
rect 303856 37924 303862 37936
rect 312630 37924 312636 37936
rect 303856 37896 312636 37924
rect 303856 37884 303862 37896
rect 312630 37884 312636 37896
rect 312688 37884 312694 37936
rect 316770 37884 316776 37936
rect 316828 37924 316834 37936
rect 327074 37924 327080 37936
rect 316828 37896 327080 37924
rect 316828 37884 316834 37896
rect 327074 37884 327080 37896
rect 327132 37884 327138 37936
rect 322934 37612 322940 37664
rect 322992 37652 322998 37664
rect 326154 37652 326160 37664
rect 322992 37624 326160 37652
rect 322992 37612 322998 37624
rect 326154 37612 326160 37624
rect 326212 37612 326218 37664
rect 297634 37204 297640 37256
rect 297692 37244 297698 37256
rect 300486 37244 300492 37256
rect 297692 37216 300492 37244
rect 297692 37204 297698 37216
rect 300486 37204 300492 37216
rect 300544 37204 300550 37256
rect 318426 37204 318432 37256
rect 318484 37244 318490 37256
rect 320818 37244 320824 37256
rect 318484 37216 320824 37244
rect 318484 37204 318490 37216
rect 320818 37204 320824 37216
rect 320876 37204 320882 37256
rect 337930 37204 337936 37256
rect 337988 37244 337994 37256
rect 340782 37244 340788 37256
rect 337988 37216 340788 37244
rect 337988 37204 337994 37216
rect 340782 37204 340788 37216
rect 340840 37204 340846 37256
rect 345658 37204 345664 37256
rect 345716 37244 345722 37256
rect 348510 37244 348516 37256
rect 345716 37216 348516 37244
rect 345716 37204 345722 37216
rect 348510 37204 348516 37216
rect 348568 37204 348574 37256
rect 318518 37136 318524 37188
rect 318576 37176 318582 37188
rect 320910 37176 320916 37188
rect 318576 37148 320916 37176
rect 318576 37136 318582 37148
rect 320910 37136 320916 37148
rect 320968 37136 320974 37188
rect 317046 37068 317052 37120
rect 317104 37108 317110 37120
rect 322750 37108 322756 37120
rect 317104 37080 322756 37108
rect 317104 37068 317110 37080
rect 322750 37068 322756 37080
rect 322808 37068 322814 37120
rect 310698 36932 310704 36984
rect 310756 36972 310762 36984
rect 316770 36972 316776 36984
rect 310756 36944 316776 36972
rect 310756 36932 310762 36944
rect 316770 36932 316776 36944
rect 316828 36932 316834 36984
rect 317322 36796 317328 36848
rect 317380 36836 317386 36848
rect 330478 36836 330484 36848
rect 317380 36808 330484 36836
rect 317380 36796 317386 36808
rect 330478 36796 330484 36808
rect 330536 36796 330542 36848
rect 283742 36728 283748 36780
rect 283800 36768 283806 36780
rect 290366 36768 290372 36780
rect 283800 36740 290372 36768
rect 283800 36728 283806 36740
rect 290366 36728 290372 36740
rect 290424 36728 290430 36780
rect 302970 36728 302976 36780
rect 303028 36768 303034 36780
rect 316862 36768 316868 36780
rect 303028 36740 316868 36768
rect 303028 36728 303034 36740
rect 316862 36728 316868 36740
rect 316920 36728 316926 36780
rect 317230 36728 317236 36780
rect 317288 36768 317294 36780
rect 330570 36768 330576 36780
rect 317288 36740 330576 36768
rect 317288 36728 317294 36740
rect 330570 36728 330576 36740
rect 330628 36728 330634 36780
rect 273898 36660 273904 36712
rect 273956 36700 273962 36712
rect 284938 36700 284944 36712
rect 273956 36672 284944 36700
rect 273956 36660 273962 36672
rect 284938 36660 284944 36672
rect 284996 36660 285002 36712
rect 302234 36660 302240 36712
rect 302292 36700 302298 36712
rect 323762 36700 323768 36712
rect 302292 36672 323768 36700
rect 302292 36660 302298 36672
rect 323762 36660 323768 36672
rect 323820 36660 323826 36712
rect 326062 36660 326068 36712
rect 326120 36700 326126 36712
rect 335998 36700 336004 36712
rect 326120 36672 336004 36700
rect 326120 36660 326126 36672
rect 335998 36660 336004 36672
rect 336056 36660 336062 36712
rect 245654 36592 245660 36644
rect 245712 36632 245718 36644
rect 273990 36632 273996 36644
rect 245712 36604 273996 36632
rect 245712 36592 245718 36604
rect 273990 36592 273996 36604
rect 274048 36592 274054 36644
rect 289722 36592 289728 36644
rect 289780 36632 289786 36644
rect 311158 36632 311164 36644
rect 289780 36604 311164 36632
rect 289780 36592 289786 36604
rect 311158 36592 311164 36604
rect 311216 36592 311222 36644
rect 323026 36592 323032 36644
rect 323084 36632 323090 36644
rect 340690 36632 340696 36644
rect 323084 36604 340696 36632
rect 323084 36592 323090 36604
rect 340690 36592 340696 36604
rect 340748 36592 340754 36644
rect 362218 36592 362224 36644
rect 362276 36632 362282 36644
rect 367738 36632 367744 36644
rect 362276 36604 367744 36632
rect 362276 36592 362282 36604
rect 367738 36592 367744 36604
rect 367796 36592 367802 36644
rect 420178 36592 420184 36644
rect 420236 36632 420242 36644
rect 429838 36632 429844 36644
rect 420236 36604 429844 36632
rect 420236 36592 420242 36604
rect 429838 36592 429844 36604
rect 429896 36592 429902 36644
rect 45554 36524 45560 36576
rect 45612 36564 45618 36576
rect 129366 36564 129372 36576
rect 45612 36536 129372 36564
rect 45612 36524 45618 36536
rect 129366 36524 129372 36536
rect 129424 36524 129430 36576
rect 176378 36524 176384 36576
rect 176436 36564 176442 36576
rect 404354 36564 404360 36576
rect 176436 36536 404360 36564
rect 176436 36524 176442 36536
rect 404354 36524 404360 36536
rect 404412 36524 404418 36576
rect 428458 36524 428464 36576
rect 428516 36564 428522 36576
rect 454862 36564 454868 36576
rect 428516 36536 454868 36564
rect 428516 36524 428522 36536
rect 454862 36524 454868 36536
rect 454920 36524 454926 36576
rect 458542 36524 458548 36576
rect 458600 36564 458606 36576
rect 463878 36564 463884 36576
rect 458600 36536 463884 36564
rect 458600 36524 458606 36536
rect 463878 36524 463884 36536
rect 463936 36524 463942 36576
rect 300762 36048 300768 36100
rect 300820 36088 300826 36100
rect 308490 36088 308496 36100
rect 300820 36060 308496 36088
rect 300820 36048 300826 36060
rect 308490 36048 308496 36060
rect 308548 36048 308554 36100
rect 377398 35300 377404 35352
rect 377456 35340 377462 35352
rect 381538 35340 381544 35352
rect 377456 35312 381544 35340
rect 377456 35300 377462 35312
rect 381538 35300 381544 35312
rect 381596 35300 381602 35352
rect 312538 35164 312544 35216
rect 312596 35204 312602 35216
rect 324314 35204 324320 35216
rect 312596 35176 324320 35204
rect 312596 35164 312602 35176
rect 324314 35164 324320 35176
rect 324372 35164 324378 35216
rect 326154 34892 326160 34944
rect 326212 34932 326218 34944
rect 333238 34932 333244 34944
rect 326212 34904 333244 34932
rect 326212 34892 326218 34904
rect 333238 34892 333244 34904
rect 333296 34892 333302 34944
rect 323670 34416 323676 34468
rect 323728 34456 323734 34468
rect 329190 34456 329196 34468
rect 323728 34428 329196 34456
rect 323728 34416 323734 34428
rect 329190 34416 329196 34428
rect 329248 34416 329254 34468
rect 340782 34416 340788 34468
rect 340840 34456 340846 34468
rect 353938 34456 353944 34468
rect 340840 34428 353944 34456
rect 340840 34416 340846 34428
rect 353938 34416 353944 34428
rect 353996 34416 354002 34468
rect 163866 34348 163872 34400
rect 163924 34388 163930 34400
rect 360194 34388 360200 34400
rect 163924 34360 360200 34388
rect 163924 34348 163930 34360
rect 360194 34348 360200 34360
rect 360252 34348 360258 34400
rect 163498 34280 163504 34332
rect 163556 34320 163562 34332
rect 416774 34320 416780 34332
rect 163556 34292 416780 34320
rect 163556 34280 163562 34292
rect 416774 34280 416780 34292
rect 416832 34280 416838 34332
rect 471238 34280 471244 34332
rect 471296 34320 471302 34332
rect 476114 34320 476120 34332
rect 471296 34292 476120 34320
rect 471296 34280 471302 34292
rect 476114 34280 476120 34292
rect 476172 34280 476178 34332
rect 163314 34212 163320 34264
rect 163372 34252 163378 34264
rect 422294 34252 422300 34264
rect 163372 34224 422300 34252
rect 163372 34212 163378 34224
rect 422294 34212 422300 34224
rect 422352 34212 422358 34264
rect 163406 34144 163412 34196
rect 163464 34184 163470 34196
rect 423674 34184 423680 34196
rect 163464 34156 423680 34184
rect 163464 34144 163470 34156
rect 423674 34144 423680 34156
rect 423732 34144 423738 34196
rect 163222 34076 163228 34128
rect 163280 34116 163286 34128
rect 427814 34116 427820 34128
rect 163280 34088 427820 34116
rect 163280 34076 163286 34088
rect 427814 34076 427820 34088
rect 427872 34076 427878 34128
rect 173158 34008 173164 34060
rect 173216 34048 173222 34060
rect 539686 34048 539692 34060
rect 173216 34020 539692 34048
rect 173216 34008 173222 34020
rect 539686 34008 539692 34020
rect 539744 34008 539750 34060
rect 173250 33940 173256 33992
rect 173308 33980 173314 33992
rect 542354 33980 542360 33992
rect 173308 33952 542360 33980
rect 173308 33940 173314 33952
rect 542354 33940 542360 33952
rect 542412 33940 542418 33992
rect 172974 33872 172980 33924
rect 173032 33912 173038 33924
rect 546494 33912 546500 33924
rect 173032 33884 546500 33912
rect 173032 33872 173038 33884
rect 546494 33872 546500 33884
rect 546552 33872 546558 33924
rect 172882 33804 172888 33856
rect 172940 33844 172946 33856
rect 552014 33844 552020 33856
rect 172940 33816 552020 33844
rect 172940 33804 172946 33816
rect 552014 33804 552020 33816
rect 552072 33804 552078 33856
rect 173066 33736 173072 33788
rect 173124 33776 173130 33788
rect 553394 33776 553400 33788
rect 173124 33748 553400 33776
rect 173124 33736 173130 33748
rect 553394 33736 553400 33748
rect 553452 33736 553458 33788
rect 337378 33124 337384 33176
rect 337436 33164 337442 33176
rect 339954 33164 339960 33176
rect 337436 33136 339960 33164
rect 337436 33124 337442 33136
rect 339954 33124 339960 33136
rect 340012 33124 340018 33176
rect 340138 33056 340144 33108
rect 340196 33096 340202 33108
rect 345934 33096 345940 33108
rect 340196 33068 345940 33096
rect 340196 33056 340202 33068
rect 345934 33056 345940 33068
rect 345992 33056 345998 33108
rect 467098 33056 467104 33108
rect 467156 33096 467162 33108
rect 472342 33096 472348 33108
rect 467156 33068 472348 33096
rect 467156 33056 467162 33068
rect 472342 33056 472348 33068
rect 472400 33056 472406 33108
rect 340690 32988 340696 33040
rect 340748 33028 340754 33040
rect 343634 33028 343640 33040
rect 340748 33000 343640 33028
rect 340748 32988 340754 33000
rect 343634 32988 343640 33000
rect 343692 32988 343698 33040
rect 3418 32784 3424 32836
rect 3476 32824 3482 32836
rect 7650 32824 7656 32836
rect 3476 32796 7656 32824
rect 3476 32784 3482 32796
rect 7650 32784 7656 32796
rect 7708 32784 7714 32836
rect 145282 32648 145288 32700
rect 145340 32688 145346 32700
rect 187694 32688 187700 32700
rect 145340 32660 187700 32688
rect 145340 32648 145346 32660
rect 187694 32648 187700 32660
rect 187752 32648 187758 32700
rect 145190 32580 145196 32632
rect 145248 32620 145254 32632
rect 194594 32620 194600 32632
rect 145248 32592 194600 32620
rect 145248 32580 145254 32592
rect 194594 32580 194600 32592
rect 194652 32580 194658 32632
rect 145374 32512 145380 32564
rect 145432 32552 145438 32564
rect 198734 32552 198740 32564
rect 145432 32524 198740 32552
rect 145432 32512 145438 32524
rect 198734 32512 198740 32524
rect 198792 32512 198798 32564
rect 369118 32512 369124 32564
rect 369176 32552 369182 32564
rect 379514 32552 379520 32564
rect 369176 32524 379520 32552
rect 369176 32512 369182 32524
rect 379514 32512 379520 32524
rect 379572 32512 379578 32564
rect 429838 32512 429844 32564
rect 429896 32552 429902 32564
rect 440878 32552 440884 32564
rect 429896 32524 440884 32552
rect 429896 32512 429902 32524
rect 440878 32512 440884 32524
rect 440936 32512 440942 32564
rect 174446 32444 174452 32496
rect 174504 32484 174510 32496
rect 556246 32484 556252 32496
rect 174504 32456 556252 32484
rect 174504 32444 174510 32456
rect 556246 32444 556252 32456
rect 556304 32444 556310 32496
rect 174354 32376 174360 32428
rect 174412 32416 174418 32428
rect 564526 32416 564532 32428
rect 174412 32388 564532 32416
rect 174412 32376 174418 32388
rect 564526 32376 564532 32388
rect 564584 32376 564590 32428
rect 336182 31832 336188 31884
rect 336240 31872 336246 31884
rect 342898 31872 342904 31884
rect 336240 31844 342904 31872
rect 336240 31832 336246 31844
rect 342898 31832 342904 31844
rect 342956 31832 342962 31884
rect 323578 31696 323584 31748
rect 323636 31736 323642 31748
rect 326338 31736 326344 31748
rect 323636 31708 326344 31736
rect 323636 31696 323642 31708
rect 326338 31696 326344 31708
rect 326396 31696 326402 31748
rect 160462 31560 160468 31612
rect 160520 31600 160526 31612
rect 382274 31600 382280 31612
rect 160520 31572 382280 31600
rect 160520 31560 160526 31572
rect 382274 31560 382280 31572
rect 382332 31560 382338 31612
rect 160554 31492 160560 31544
rect 160612 31532 160618 31544
rect 389174 31532 389180 31544
rect 160612 31504 389180 31532
rect 160612 31492 160618 31504
rect 389174 31492 389180 31504
rect 389232 31492 389238 31544
rect 163038 31424 163044 31476
rect 163096 31464 163102 31476
rect 423766 31464 423772 31476
rect 163096 31436 423772 31464
rect 163096 31424 163102 31436
rect 423766 31424 423772 31436
rect 423824 31424 423830 31476
rect 163130 31356 163136 31408
rect 163188 31396 163194 31408
rect 426434 31396 426440 31408
rect 163188 31368 426440 31396
rect 163188 31356 163194 31368
rect 426434 31356 426440 31368
rect 426492 31356 426498 31408
rect 454862 31356 454868 31408
rect 454920 31396 454926 31408
rect 458818 31396 458824 31408
rect 454920 31368 458824 31396
rect 454920 31356 454926 31368
rect 458818 31356 458824 31368
rect 458876 31356 458882 31408
rect 164510 31288 164516 31340
rect 164568 31328 164574 31340
rect 438854 31328 438860 31340
rect 164568 31300 438860 31328
rect 164568 31288 164574 31300
rect 438854 31288 438860 31300
rect 438912 31288 438918 31340
rect 463878 31288 463884 31340
rect 463936 31328 463942 31340
rect 473354 31328 473360 31340
rect 463936 31300 473360 31328
rect 463936 31288 463942 31300
rect 473354 31288 473360 31300
rect 473412 31288 473418 31340
rect 172514 31220 172520 31272
rect 172572 31260 172578 31272
rect 540974 31260 540980 31272
rect 172572 31232 540980 31260
rect 172572 31220 172578 31232
rect 540974 31220 540980 31232
rect 541032 31220 541038 31272
rect 172606 31152 172612 31204
rect 172664 31192 172670 31204
rect 545114 31192 545120 31204
rect 172664 31164 545120 31192
rect 172664 31152 172670 31164
rect 545114 31152 545120 31164
rect 545172 31152 545178 31204
rect 172698 31084 172704 31136
rect 172756 31124 172762 31136
rect 547966 31124 547972 31136
rect 172756 31096 547972 31124
rect 172756 31084 172762 31096
rect 547966 31084 547972 31096
rect 548024 31084 548030 31136
rect 172790 31016 172796 31068
rect 172848 31056 172854 31068
rect 550634 31056 550640 31068
rect 172848 31028 550640 31056
rect 172848 31016 172854 31028
rect 550634 31016 550640 31028
rect 550692 31016 550698 31068
rect 327074 30948 327080 31000
rect 327132 30988 327138 31000
rect 330662 30988 330668 31000
rect 327132 30960 330668 30988
rect 327132 30948 327138 30960
rect 330662 30948 330668 30960
rect 330720 30948 330726 31000
rect 300486 30268 300492 30320
rect 300544 30308 300550 30320
rect 302234 30308 302240 30320
rect 300544 30280 302240 30308
rect 300544 30268 300550 30280
rect 302234 30268 302240 30280
rect 302292 30268 302298 30320
rect 325050 30268 325056 30320
rect 325108 30308 325114 30320
rect 327902 30308 327908 30320
rect 325108 30280 327908 30308
rect 325108 30268 325114 30280
rect 327902 30268 327908 30280
rect 327960 30268 327966 30320
rect 339954 30268 339960 30320
rect 340012 30308 340018 30320
rect 345014 30308 345020 30320
rect 340012 30280 345020 30308
rect 340012 30268 340018 30280
rect 345014 30268 345020 30280
rect 345072 30268 345078 30320
rect 343634 30200 343640 30252
rect 343692 30240 343698 30252
rect 347038 30240 347044 30252
rect 343692 30212 347044 30240
rect 343692 30200 343698 30212
rect 347038 30200 347044 30212
rect 347096 30200 347102 30252
rect 290366 29656 290372 29708
rect 290424 29696 290430 29708
rect 309778 29696 309784 29708
rect 290424 29668 309784 29696
rect 290424 29656 290430 29668
rect 309778 29656 309784 29668
rect 309836 29656 309842 29708
rect 322750 29656 322756 29708
rect 322808 29696 322814 29708
rect 344462 29696 344468 29708
rect 322808 29668 344468 29696
rect 322808 29656 322814 29668
rect 344462 29656 344468 29668
rect 344520 29656 344526 29708
rect 472342 29656 472348 29708
rect 472400 29696 472406 29708
rect 477494 29696 477500 29708
rect 472400 29668 477500 29696
rect 472400 29656 472406 29668
rect 477494 29656 477500 29668
rect 477552 29656 477558 29708
rect 168742 29588 168748 29640
rect 168800 29628 168806 29640
rect 490006 29628 490012 29640
rect 168800 29600 490012 29628
rect 168800 29588 168806 29600
rect 490006 29588 490012 29600
rect 490064 29588 490070 29640
rect 154022 28908 154028 28960
rect 154080 28948 154086 28960
rect 289814 28948 289820 28960
rect 154080 28920 289820 28948
rect 154080 28908 154086 28920
rect 289814 28908 289820 28920
rect 289872 28908 289878 28960
rect 308490 28908 308496 28960
rect 308548 28948 308554 28960
rect 316586 28948 316592 28960
rect 308548 28920 316592 28948
rect 308548 28908 308554 28920
rect 316586 28908 316592 28920
rect 316644 28908 316650 28960
rect 316862 28908 316868 28960
rect 316920 28948 316926 28960
rect 319622 28948 319628 28960
rect 316920 28920 319628 28948
rect 316920 28908 316926 28920
rect 319622 28908 319628 28920
rect 319680 28908 319686 28960
rect 336090 28908 336096 28960
rect 336148 28948 336154 28960
rect 341058 28948 341064 28960
rect 336148 28920 341064 28948
rect 336148 28908 336154 28920
rect 341058 28908 341064 28920
rect 341116 28908 341122 28960
rect 347130 28908 347136 28960
rect 347188 28948 347194 28960
rect 352558 28948 352564 28960
rect 347188 28920 352564 28948
rect 347188 28908 347194 28920
rect 352558 28908 352564 28920
rect 352616 28908 352622 28960
rect 379514 28908 379520 28960
rect 379572 28948 379578 28960
rect 382918 28948 382924 28960
rect 379572 28920 382924 28948
rect 379572 28908 379578 28920
rect 382918 28908 382924 28920
rect 382976 28908 382982 28960
rect 166626 28840 166632 28892
rect 166684 28880 166690 28892
rect 375374 28880 375380 28892
rect 166684 28852 375380 28880
rect 166684 28840 166690 28852
rect 375374 28840 375380 28852
rect 375432 28840 375438 28892
rect 166534 28772 166540 28824
rect 166592 28812 166598 28824
rect 397454 28812 397460 28824
rect 166592 28784 397460 28812
rect 166592 28772 166598 28784
rect 397454 28772 397460 28784
rect 397512 28772 397518 28824
rect 162026 28704 162032 28756
rect 162084 28744 162090 28756
rect 407114 28744 407120 28756
rect 162084 28716 407120 28744
rect 162084 28704 162090 28716
rect 407114 28704 407120 28716
rect 407172 28704 407178 28756
rect 162946 28636 162952 28688
rect 163004 28676 163010 28688
rect 415486 28676 415492 28688
rect 163004 28648 415492 28676
rect 163004 28636 163010 28648
rect 415486 28636 415492 28648
rect 415544 28636 415550 28688
rect 166166 28568 166172 28620
rect 166224 28608 166230 28620
rect 449894 28608 449900 28620
rect 166224 28580 449900 28608
rect 166224 28568 166230 28580
rect 449894 28568 449900 28580
rect 449952 28568 449958 28620
rect 165982 28500 165988 28552
rect 166040 28540 166046 28552
rect 452654 28540 452660 28552
rect 166040 28512 452660 28540
rect 166040 28500 166046 28512
rect 452654 28500 452660 28512
rect 452712 28500 452718 28552
rect 166074 28432 166080 28484
rect 166132 28472 166138 28484
rect 456886 28472 456892 28484
rect 166132 28444 456892 28472
rect 166132 28432 166138 28444
rect 456886 28432 456892 28444
rect 456944 28432 456950 28484
rect 166258 28364 166264 28416
rect 166316 28404 166322 28416
rect 459554 28404 459560 28416
rect 166316 28376 459560 28404
rect 166316 28364 166322 28376
rect 459554 28364 459560 28376
rect 459612 28364 459618 28416
rect 171686 28296 171692 28348
rect 171744 28336 171750 28348
rect 521654 28336 521660 28348
rect 171744 28308 521660 28336
rect 171744 28296 171750 28308
rect 521654 28296 521660 28308
rect 521712 28296 521718 28348
rect 171594 28228 171600 28280
rect 171652 28268 171658 28280
rect 524414 28268 524420 28280
rect 171652 28240 524420 28268
rect 171652 28228 171658 28240
rect 524414 28228 524420 28240
rect 524472 28228 524478 28280
rect 146938 28160 146944 28212
rect 146996 28200 147002 28212
rect 209774 28200 209780 28212
rect 146996 28172 209780 28200
rect 146996 28160 147002 28172
rect 209774 28160 209780 28172
rect 209832 28160 209838 28212
rect 316586 28160 316592 28212
rect 316644 28200 316650 28212
rect 318058 28200 318064 28212
rect 316644 28172 318064 28200
rect 316644 28160 316650 28172
rect 318058 28160 318064 28172
rect 318116 28160 318122 28212
rect 345934 28160 345940 28212
rect 345992 28200 345998 28212
rect 353294 28200 353300 28212
rect 345992 28172 353300 28200
rect 345992 28160 345998 28172
rect 353294 28160 353300 28172
rect 353352 28160 353358 28212
rect 146846 28092 146852 28144
rect 146904 28132 146910 28144
rect 205634 28132 205640 28144
rect 146904 28104 205640 28132
rect 146904 28092 146910 28104
rect 205634 28092 205640 28104
rect 205692 28092 205698 28144
rect 146754 28024 146760 28076
rect 146812 28064 146818 28076
rect 201494 28064 201500 28076
rect 146812 28036 201500 28064
rect 146812 28024 146818 28036
rect 201494 28024 201500 28036
rect 201552 28024 201558 28076
rect 324958 27616 324964 27668
rect 325016 27656 325022 27668
rect 327074 27656 327080 27668
rect 325016 27628 327080 27656
rect 325016 27616 325022 27628
rect 327074 27616 327080 27628
rect 327132 27616 327138 27668
rect 307018 27548 307024 27600
rect 307076 27588 307082 27600
rect 312170 27588 312176 27600
rect 307076 27560 312176 27588
rect 307076 27548 307082 27560
rect 312170 27548 312176 27560
rect 312228 27548 312234 27600
rect 348510 27548 348516 27600
rect 348568 27588 348574 27600
rect 352650 27588 352656 27600
rect 348568 27560 352656 27588
rect 348568 27548 348574 27560
rect 352650 27548 352656 27560
rect 352708 27548 352714 27600
rect 312630 27004 312636 27056
rect 312688 27044 312694 27056
rect 320082 27044 320088 27056
rect 312688 27016 320088 27044
rect 312688 27004 312694 27016
rect 320082 27004 320088 27016
rect 320140 27004 320146 27056
rect 323762 27004 323768 27056
rect 323820 27044 323826 27056
rect 329098 27044 329104 27056
rect 323820 27016 329104 27044
rect 323820 27004 323826 27016
rect 329098 27004 329104 27016
rect 329156 27004 329162 27056
rect 145098 26936 145104 26988
rect 145156 26976 145162 26988
rect 193306 26976 193312 26988
rect 145156 26948 193312 26976
rect 145156 26936 145162 26948
rect 193306 26936 193312 26948
rect 193364 26936 193370 26988
rect 300118 26936 300124 26988
rect 300176 26976 300182 26988
rect 321186 26976 321192 26988
rect 300176 26948 321192 26976
rect 300176 26936 300182 26948
rect 321186 26936 321192 26948
rect 321244 26936 321250 26988
rect 324314 26936 324320 26988
rect 324372 26976 324378 26988
rect 334618 26976 334624 26988
rect 324372 26948 334624 26976
rect 324372 26936 324378 26948
rect 334618 26936 334624 26948
rect 334676 26936 334682 26988
rect 160370 26868 160376 26920
rect 160428 26908 160434 26920
rect 385034 26908 385040 26920
rect 160428 26880 385040 26908
rect 160428 26868 160434 26880
rect 385034 26868 385040 26880
rect 385092 26868 385098 26920
rect 439498 26868 439504 26920
rect 439556 26908 439562 26920
rect 446398 26908 446404 26920
rect 439556 26880 446404 26908
rect 439556 26868 439562 26880
rect 446398 26868 446404 26880
rect 446456 26868 446462 26920
rect 464338 26868 464344 26920
rect 464396 26908 464402 26920
rect 493318 26908 493324 26920
rect 464396 26880 493324 26908
rect 464396 26868 464402 26880
rect 493318 26868 493324 26880
rect 493376 26868 493382 26920
rect 302234 26324 302240 26376
rect 302292 26364 302298 26376
rect 306374 26364 306380 26376
rect 302292 26336 306380 26364
rect 302292 26324 302298 26336
rect 306374 26324 306380 26336
rect 306432 26324 306438 26376
rect 283558 26120 283564 26172
rect 283616 26160 283622 26172
rect 292758 26160 292764 26172
rect 283616 26132 292764 26160
rect 283616 26120 283622 26132
rect 292758 26120 292764 26132
rect 292816 26120 292822 26172
rect 145006 26052 145012 26104
rect 145064 26092 145070 26104
rect 186314 26092 186320 26104
rect 145064 26064 186320 26092
rect 145064 26052 145070 26064
rect 186314 26052 186320 26064
rect 186372 26052 186378 26104
rect 283650 26052 283656 26104
rect 283708 26092 283714 26104
rect 294046 26092 294052 26104
rect 283708 26064 294052 26092
rect 283708 26052 283714 26064
rect 294046 26052 294052 26064
rect 294104 26052 294110 26104
rect 363598 26052 363604 26104
rect 363656 26092 363662 26104
rect 367554 26092 367560 26104
rect 363656 26064 367560 26092
rect 363656 26052 363662 26064
rect 367554 26052 367560 26064
rect 367612 26052 367618 26104
rect 152734 25984 152740 26036
rect 152792 26024 152798 26036
rect 253934 26024 253940 26036
rect 152792 25996 253940 26024
rect 152792 25984 152798 25996
rect 253934 25984 253940 25996
rect 253992 25984 253998 26036
rect 280798 25984 280804 26036
rect 280856 26024 280862 26036
rect 294138 26024 294144 26036
rect 280856 25996 294144 26024
rect 280856 25984 280862 25996
rect 294138 25984 294144 25996
rect 294196 25984 294202 26036
rect 315298 25984 315304 26036
rect 315356 26024 315362 26036
rect 320174 26024 320180 26036
rect 315356 25996 320180 26024
rect 315356 25984 315362 25996
rect 320174 25984 320180 25996
rect 320232 25984 320238 26036
rect 321094 25984 321100 26036
rect 321152 26024 321158 26036
rect 329006 26024 329012 26036
rect 321152 25996 329012 26024
rect 321152 25984 321158 25996
rect 329006 25984 329012 25996
rect 329064 25984 329070 26036
rect 333238 25984 333244 26036
rect 333296 26024 333302 26036
rect 343634 26024 343640 26036
rect 333296 25996 343640 26024
rect 333296 25984 333302 25996
rect 343634 25984 343640 25996
rect 343692 25984 343698 26036
rect 349798 25984 349804 26036
rect 349856 26024 349862 26036
rect 364978 26024 364984 26036
rect 349856 25996 364984 26024
rect 349856 25984 349862 25996
rect 364978 25984 364984 25996
rect 365036 25984 365042 26036
rect 162578 25916 162584 25968
rect 162636 25956 162642 25968
rect 368474 25956 368480 25968
rect 162636 25928 368480 25956
rect 162636 25916 162642 25928
rect 368474 25916 368480 25928
rect 368532 25916 368538 25968
rect 162486 25848 162492 25900
rect 162544 25888 162550 25900
rect 390554 25888 390560 25900
rect 162544 25860 390560 25888
rect 162544 25848 162550 25860
rect 390554 25848 390560 25860
rect 390612 25848 390618 25900
rect 170214 25780 170220 25832
rect 170272 25820 170278 25832
rect 506474 25820 506480 25832
rect 170272 25792 506480 25820
rect 170272 25780 170278 25792
rect 506474 25780 506480 25792
rect 506532 25780 506538 25832
rect 171502 25712 171508 25764
rect 171560 25752 171566 25764
rect 528554 25752 528560 25764
rect 171560 25724 528560 25752
rect 171560 25712 171566 25724
rect 528554 25712 528560 25724
rect 528612 25712 528618 25764
rect 174170 25644 174176 25696
rect 174228 25684 174234 25696
rect 558914 25684 558920 25696
rect 174228 25656 558920 25684
rect 174228 25644 174234 25656
rect 558914 25644 558920 25656
rect 558972 25644 558978 25696
rect 174078 25576 174084 25628
rect 174136 25616 174142 25628
rect 563054 25616 563060 25628
rect 174136 25588 563060 25616
rect 174136 25576 174142 25588
rect 563054 25576 563060 25588
rect 563112 25576 563118 25628
rect 174262 25508 174268 25560
rect 174320 25548 174326 25560
rect 565814 25548 565820 25560
rect 174320 25520 565820 25548
rect 174320 25508 174326 25520
rect 565814 25508 565820 25520
rect 565872 25508 565878 25560
rect 302878 24828 302884 24880
rect 302936 24868 302942 24880
rect 307110 24868 307116 24880
rect 302936 24840 307116 24868
rect 302936 24828 302942 24840
rect 307110 24828 307116 24840
rect 307168 24828 307174 24880
rect 321002 24828 321008 24880
rect 321060 24868 321066 24880
rect 323578 24868 323584 24880
rect 321060 24840 323584 24868
rect 321060 24828 321066 24840
rect 323578 24828 323584 24840
rect 323636 24828 323642 24880
rect 291838 24556 291844 24608
rect 291896 24596 291902 24608
rect 294322 24596 294328 24608
rect 291896 24568 294328 24596
rect 291896 24556 291902 24568
rect 294322 24556 294328 24568
rect 294380 24556 294386 24608
rect 316770 24420 316776 24472
rect 316828 24460 316834 24472
rect 319530 24460 319536 24472
rect 316828 24432 319536 24460
rect 316828 24420 316834 24432
rect 319530 24420 319536 24432
rect 319588 24420 319594 24472
rect 440878 24284 440884 24336
rect 440936 24324 440942 24336
rect 443730 24324 443736 24336
rect 440936 24296 443736 24324
rect 440936 24284 440942 24296
rect 443730 24284 443736 24296
rect 443788 24284 443794 24336
rect 292022 24216 292028 24268
rect 292080 24256 292086 24268
rect 300670 24256 300676 24268
rect 292080 24228 300676 24256
rect 292080 24216 292086 24228
rect 300670 24216 300676 24228
rect 300728 24216 300734 24268
rect 273990 24148 273996 24200
rect 274048 24188 274054 24200
rect 292666 24188 292672 24200
rect 274048 24160 292672 24188
rect 274048 24148 274054 24160
rect 292666 24148 292672 24160
rect 292724 24148 292730 24200
rect 320082 24148 320088 24200
rect 320140 24188 320146 24200
rect 324958 24188 324964 24200
rect 320140 24160 324964 24188
rect 320140 24148 320146 24160
rect 324958 24148 324964 24160
rect 325016 24148 325022 24200
rect 327902 24148 327908 24200
rect 327960 24188 327966 24200
rect 344370 24188 344376 24200
rect 327960 24160 344376 24188
rect 327960 24148 327966 24160
rect 344370 24148 344376 24160
rect 344428 24148 344434 24200
rect 2958 24080 2964 24132
rect 3016 24120 3022 24132
rect 189166 24120 189172 24132
rect 3016 24092 189172 24120
rect 3016 24080 3022 24092
rect 189166 24080 189172 24092
rect 189224 24080 189230 24132
rect 284938 24080 284944 24132
rect 284996 24120 285002 24132
rect 304442 24120 304448 24132
rect 284996 24092 304448 24120
rect 284996 24080 285002 24092
rect 304442 24080 304448 24092
rect 304500 24080 304506 24132
rect 326338 24080 326344 24132
rect 326396 24120 326402 24132
rect 342254 24120 342260 24132
rect 326396 24092 342260 24120
rect 326396 24080 326402 24092
rect 342254 24080 342260 24092
rect 342312 24080 342318 24132
rect 344462 24080 344468 24132
rect 344520 24120 344526 24132
rect 349890 24120 349896 24132
rect 344520 24092 349896 24120
rect 344520 24080 344526 24092
rect 349890 24080 349896 24092
rect 349948 24080 349954 24132
rect 353294 24080 353300 24132
rect 353352 24120 353358 24132
rect 359274 24120 359280 24132
rect 353352 24092 359280 24120
rect 353352 24080 353358 24092
rect 359274 24080 359280 24092
rect 359332 24080 359338 24132
rect 141234 23400 141240 23452
rect 141292 23440 141298 23452
rect 142154 23440 142160 23452
rect 141292 23412 142160 23440
rect 141292 23400 141298 23412
rect 142154 23400 142160 23412
rect 142212 23400 142218 23452
rect 146662 23400 146668 23452
rect 146720 23440 146726 23452
rect 204254 23440 204260 23452
rect 146720 23412 204260 23440
rect 146720 23400 146726 23412
rect 204254 23400 204260 23412
rect 204312 23400 204318 23452
rect 381538 23400 381544 23452
rect 381596 23440 381602 23452
rect 384298 23440 384304 23452
rect 381596 23412 384304 23440
rect 381596 23400 381602 23412
rect 384298 23400 384304 23412
rect 384356 23400 384362 23452
rect 146478 23332 146484 23384
rect 146536 23372 146542 23384
rect 208394 23372 208400 23384
rect 146536 23344 208400 23372
rect 146536 23332 146542 23344
rect 208394 23332 208400 23344
rect 208452 23332 208458 23384
rect 146570 23264 146576 23316
rect 146628 23304 146634 23316
rect 211154 23304 211160 23316
rect 146628 23276 211160 23304
rect 146628 23264 146634 23276
rect 211154 23264 211160 23276
rect 211212 23264 211218 23316
rect 272518 23264 272524 23316
rect 272576 23304 272582 23316
rect 275002 23304 275008 23316
rect 272576 23276 275008 23304
rect 272576 23264 272582 23276
rect 275002 23264 275008 23276
rect 275060 23264 275066 23316
rect 309778 23264 309784 23316
rect 309836 23304 309842 23316
rect 312906 23304 312912 23316
rect 309836 23276 312912 23304
rect 309836 23264 309842 23276
rect 312906 23264 312912 23276
rect 312964 23264 312970 23316
rect 152458 23196 152464 23248
rect 152516 23236 152522 23248
rect 273254 23236 273260 23248
rect 152516 23208 273260 23236
rect 152516 23196 152522 23208
rect 273254 23196 273260 23208
rect 273312 23196 273318 23248
rect 308398 23196 308404 23248
rect 308456 23236 308462 23248
rect 313274 23236 313280 23248
rect 308456 23208 313280 23236
rect 308456 23196 308462 23208
rect 313274 23196 313280 23208
rect 313332 23196 313338 23248
rect 152366 23128 152372 23180
rect 152424 23168 152430 23180
rect 280154 23168 280160 23180
rect 152424 23140 280160 23168
rect 152424 23128 152430 23140
rect 280154 23128 280160 23140
rect 280212 23128 280218 23180
rect 142614 23060 142620 23112
rect 142672 23100 142678 23112
rect 149054 23100 149060 23112
rect 142672 23072 149060 23100
rect 142672 23060 142678 23072
rect 149054 23060 149060 23072
rect 149112 23060 149118 23112
rect 153746 23060 153752 23112
rect 153804 23100 153810 23112
rect 291194 23100 291200 23112
rect 153804 23072 291200 23100
rect 153804 23060 153810 23072
rect 291194 23060 291200 23072
rect 291252 23060 291258 23112
rect 141326 22992 141332 23044
rect 141384 23032 141390 23044
rect 145006 23032 145012 23044
rect 141384 23004 145012 23032
rect 141384 22992 141390 23004
rect 145006 22992 145012 23004
rect 145064 22992 145070 23044
rect 153930 22992 153936 23044
rect 153988 23032 153994 23044
rect 293954 23032 293960 23044
rect 153988 23004 293960 23032
rect 153988 22992 153994 23004
rect 293954 22992 293960 23004
rect 294012 22992 294018 23044
rect 294598 22992 294604 23044
rect 294656 23032 294662 23044
rect 305638 23032 305644 23044
rect 294656 23004 305644 23032
rect 294656 22992 294662 23004
rect 305638 22992 305644 23004
rect 305696 22992 305702 23044
rect 153838 22924 153844 22976
rect 153896 22964 153902 22976
rect 300854 22964 300860 22976
rect 153896 22936 300860 22964
rect 153896 22924 153902 22936
rect 300854 22924 300860 22936
rect 300912 22924 300918 22976
rect 3418 22856 3424 22908
rect 3476 22896 3482 22908
rect 178126 22896 178132 22908
rect 3476 22868 178132 22896
rect 3476 22856 3482 22868
rect 178126 22856 178132 22868
rect 178184 22856 178190 22908
rect 291930 22856 291936 22908
rect 291988 22896 291994 22908
rect 307018 22896 307024 22908
rect 291988 22868 307024 22896
rect 291988 22856 291994 22868
rect 307018 22856 307024 22868
rect 307076 22856 307082 22908
rect 129642 22788 129648 22840
rect 129700 22828 129706 22840
rect 304994 22828 305000 22840
rect 129700 22800 305000 22828
rect 129700 22788 129706 22800
rect 304994 22788 305000 22800
rect 305052 22788 305058 22840
rect 306374 22788 306380 22840
rect 306432 22828 306438 22840
rect 340046 22828 340052 22840
rect 306432 22800 340052 22828
rect 306432 22788 306438 22800
rect 340046 22788 340052 22800
rect 340104 22788 340110 22840
rect 341058 22788 341064 22840
rect 341116 22828 341122 22840
rect 358078 22828 358084 22840
rect 341116 22800 358084 22828
rect 341116 22788 341122 22800
rect 358078 22788 358084 22800
rect 358136 22788 358142 22840
rect 120718 22720 120724 22772
rect 120776 22760 120782 22772
rect 580258 22760 580264 22772
rect 120776 22732 580264 22760
rect 120776 22720 120782 22732
rect 580258 22720 580264 22732
rect 580316 22720 580322 22772
rect 329006 22652 329012 22704
rect 329064 22692 329070 22704
rect 334802 22692 334808 22704
rect 329064 22664 334808 22692
rect 329064 22652 329070 22664
rect 334802 22652 334808 22664
rect 334860 22652 334866 22704
rect 312170 22312 312176 22364
rect 312228 22352 312234 22364
rect 315298 22352 315304 22364
rect 312228 22324 315304 22352
rect 312228 22312 312234 22324
rect 315298 22312 315304 22324
rect 315356 22312 315362 22364
rect 294322 22040 294328 22092
rect 294380 22080 294386 22092
rect 298002 22080 298008 22092
rect 294380 22052 298008 22080
rect 294380 22040 294386 22052
rect 298002 22040 298008 22052
rect 298060 22040 298066 22092
rect 352650 22040 352656 22092
rect 352708 22080 352714 22092
rect 357158 22080 357164 22092
rect 352708 22052 357164 22080
rect 352708 22040 352714 22052
rect 357158 22040 357164 22052
rect 357216 22040 357222 22092
rect 446398 22040 446404 22092
rect 446456 22080 446462 22092
rect 448882 22080 448888 22092
rect 446456 22052 448888 22080
rect 446456 22040 446462 22052
rect 448882 22040 448888 22052
rect 448940 22040 448946 22092
rect 329190 21700 329196 21752
rect 329248 21740 329254 21752
rect 341518 21740 341524 21752
rect 329248 21712 341524 21740
rect 329248 21700 329254 21712
rect 341518 21700 341524 21712
rect 341576 21700 341582 21752
rect 327074 21632 327080 21684
rect 327132 21672 327138 21684
rect 340138 21672 340144 21684
rect 327132 21644 340144 21672
rect 327132 21632 327138 21644
rect 340138 21632 340144 21644
rect 340196 21632 340202 21684
rect 344278 21632 344284 21684
rect 344336 21672 344342 21684
rect 352650 21672 352656 21684
rect 344336 21644 352656 21672
rect 344336 21632 344342 21644
rect 352650 21632 352656 21644
rect 352708 21632 352714 21684
rect 177666 21564 177672 21616
rect 177724 21604 177730 21616
rect 418154 21604 418160 21616
rect 177724 21576 418160 21604
rect 177724 21564 177730 21576
rect 418154 21564 418160 21576
rect 418212 21564 418218 21616
rect 169938 21496 169944 21548
rect 169996 21536 170002 21548
rect 506566 21536 506572 21548
rect 169996 21508 506572 21536
rect 169996 21496 170002 21508
rect 506566 21496 506572 21508
rect 506624 21496 506630 21548
rect 170122 21428 170128 21480
rect 170180 21468 170186 21480
rect 509234 21468 509240 21480
rect 170180 21440 509240 21468
rect 170180 21428 170186 21440
rect 509234 21428 509240 21440
rect 509292 21428 509298 21480
rect 170030 21360 170036 21412
rect 170088 21400 170094 21412
rect 513374 21400 513380 21412
rect 170088 21372 513380 21400
rect 170088 21360 170094 21372
rect 513374 21360 513380 21372
rect 513432 21360 513438 21412
rect 150894 20612 150900 20664
rect 150952 20652 150958 20664
rect 255314 20652 255320 20664
rect 150952 20624 255320 20652
rect 150952 20612 150958 20624
rect 255314 20612 255320 20624
rect 255372 20612 255378 20664
rect 300670 20612 300676 20664
rect 300728 20652 300734 20664
rect 308490 20652 308496 20664
rect 300728 20624 308496 20652
rect 300728 20612 300734 20624
rect 308490 20612 308496 20624
rect 308548 20612 308554 20664
rect 347038 20612 347044 20664
rect 347096 20652 347102 20664
rect 349798 20652 349804 20664
rect 347096 20624 349804 20652
rect 347096 20612 347102 20624
rect 349798 20612 349804 20624
rect 349856 20612 349862 20664
rect 349890 20612 349896 20664
rect 349948 20652 349954 20664
rect 355594 20652 355600 20664
rect 349948 20624 355600 20652
rect 349948 20612 349954 20624
rect 355594 20612 355600 20624
rect 355652 20612 355658 20664
rect 359274 20612 359280 20664
rect 359332 20652 359338 20664
rect 365070 20652 365076 20664
rect 359332 20624 365076 20652
rect 359332 20612 359338 20624
rect 365070 20612 365076 20624
rect 365128 20612 365134 20664
rect 367554 20612 367560 20664
rect 367612 20652 367618 20664
rect 371234 20652 371240 20664
rect 367612 20624 371240 20652
rect 367612 20612 367618 20624
rect 371234 20612 371240 20624
rect 371292 20612 371298 20664
rect 526438 20612 526444 20664
rect 526496 20652 526502 20664
rect 579982 20652 579988 20664
rect 526496 20624 579988 20652
rect 526496 20612 526502 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 150986 20544 150992 20596
rect 151044 20584 151050 20596
rect 259546 20584 259552 20596
rect 151044 20556 259552 20584
rect 151044 20544 151050 20556
rect 259546 20544 259552 20556
rect 259604 20544 259610 20596
rect 151078 20476 151084 20528
rect 151136 20516 151142 20528
rect 262214 20516 262220 20528
rect 151136 20488 262220 20516
rect 151136 20476 151142 20488
rect 262214 20476 262220 20488
rect 262272 20476 262278 20528
rect 151170 20408 151176 20460
rect 151228 20448 151234 20460
rect 269114 20448 269120 20460
rect 151228 20420 269120 20448
rect 151228 20408 151234 20420
rect 269114 20408 269120 20420
rect 269172 20408 269178 20460
rect 275002 20408 275008 20460
rect 275060 20448 275066 20460
rect 288342 20448 288348 20460
rect 275060 20420 288348 20448
rect 275060 20408 275066 20420
rect 288342 20408 288348 20420
rect 288400 20408 288406 20460
rect 292666 20408 292672 20460
rect 292724 20448 292730 20460
rect 300118 20448 300124 20460
rect 292724 20420 300124 20448
rect 292724 20408 292730 20420
rect 300118 20408 300124 20420
rect 300176 20408 300182 20460
rect 152274 20340 152280 20392
rect 152332 20380 152338 20392
rect 276014 20380 276020 20392
rect 152332 20352 276020 20380
rect 152332 20340 152338 20352
rect 276014 20340 276020 20352
rect 276072 20340 276078 20392
rect 292758 20340 292764 20392
rect 292816 20380 292822 20392
rect 307202 20380 307208 20392
rect 292816 20352 307208 20380
rect 292816 20340 292822 20352
rect 307202 20340 307208 20352
rect 307260 20340 307266 20392
rect 153654 20272 153660 20324
rect 153712 20312 153718 20324
rect 298094 20312 298100 20324
rect 153712 20284 298100 20312
rect 153712 20272 153718 20284
rect 298094 20272 298100 20284
rect 298152 20272 298158 20324
rect 312906 20272 312912 20324
rect 312964 20312 312970 20324
rect 327074 20312 327080 20324
rect 312964 20284 327080 20312
rect 312964 20272 312970 20284
rect 327074 20272 327080 20284
rect 327132 20272 327138 20324
rect 161934 20204 161940 20256
rect 161992 20244 161998 20256
rect 402974 20244 402980 20256
rect 161992 20216 402980 20244
rect 161992 20204 161998 20216
rect 402974 20204 402980 20216
rect 403032 20204 403038 20256
rect 170950 20136 170956 20188
rect 171008 20176 171014 20188
rect 488534 20176 488540 20188
rect 171008 20148 488540 20176
rect 171008 20136 171014 20148
rect 488534 20136 488540 20148
rect 488592 20136 488598 20188
rect 168650 20068 168656 20120
rect 168708 20108 168714 20120
rect 495434 20108 495440 20120
rect 168708 20080 495440 20108
rect 168708 20068 168714 20080
rect 495434 20068 495440 20080
rect 495492 20068 495498 20120
rect 168558 20000 168564 20052
rect 168616 20040 168622 20052
rect 498286 20040 498292 20052
rect 168616 20012 498292 20040
rect 168616 20000 168622 20012
rect 498286 20000 498292 20012
rect 498344 20000 498350 20052
rect 120074 19932 120080 19984
rect 120132 19972 120138 19984
rect 139670 19972 139676 19984
rect 120132 19944 139676 19972
rect 120132 19932 120138 19944
rect 139670 19932 139676 19944
rect 139728 19932 139734 19984
rect 171410 19932 171416 19984
rect 171468 19972 171474 19984
rect 531406 19972 531412 19984
rect 171468 19944 531412 19972
rect 171468 19932 171474 19944
rect 531406 19932 531412 19944
rect 531464 19932 531470 19984
rect 149698 19864 149704 19916
rect 149756 19904 149762 19916
rect 237374 19904 237380 19916
rect 149756 19876 237380 19904
rect 149756 19864 149762 19876
rect 237374 19864 237380 19876
rect 237432 19864 237438 19916
rect 330662 19252 330668 19304
rect 330720 19292 330726 19304
rect 334710 19292 334716 19304
rect 330720 19264 334716 19292
rect 330720 19252 330726 19264
rect 334710 19252 334716 19264
rect 334768 19252 334774 19304
rect 330570 18776 330576 18828
rect 330628 18816 330634 18828
rect 338758 18816 338764 18828
rect 330628 18788 338764 18816
rect 330628 18776 330634 18788
rect 338758 18776 338764 18788
rect 338816 18776 338822 18828
rect 448882 18776 448888 18828
rect 448940 18816 448946 18828
rect 452746 18816 452752 18828
rect 448940 18788 452752 18816
rect 448940 18776 448946 18788
rect 452746 18776 452752 18788
rect 452804 18776 452810 18828
rect 294046 18708 294052 18760
rect 294104 18748 294110 18760
rect 304350 18748 304356 18760
rect 294104 18720 304356 18748
rect 294104 18708 294110 18720
rect 304350 18708 304356 18720
rect 304408 18708 304414 18760
rect 146202 18640 146208 18692
rect 146260 18680 146266 18692
rect 218054 18680 218060 18692
rect 146260 18652 218060 18680
rect 146260 18640 146266 18652
rect 218054 18640 218060 18652
rect 218112 18640 218118 18692
rect 298002 18640 298008 18692
rect 298060 18680 298066 18692
rect 312538 18680 312544 18692
rect 298060 18652 312544 18680
rect 298060 18640 298066 18652
rect 312538 18640 312544 18652
rect 312596 18640 312602 18692
rect 330478 18640 330484 18692
rect 330536 18680 330542 18692
rect 339310 18680 339316 18692
rect 330536 18652 339316 18680
rect 330536 18640 330542 18652
rect 339310 18640 339316 18652
rect 339368 18640 339374 18692
rect 340138 18640 340144 18692
rect 340196 18680 340202 18692
rect 349154 18680 349160 18692
rect 340196 18652 349160 18680
rect 340196 18640 340202 18652
rect 349154 18640 349160 18652
rect 349212 18640 349218 18692
rect 357158 18640 357164 18692
rect 357216 18680 357222 18692
rect 369118 18680 369124 18692
rect 357216 18652 369124 18680
rect 357216 18640 357222 18652
rect 369118 18640 369124 18652
rect 369176 18640 369182 18692
rect 173986 18572 173992 18624
rect 174044 18612 174050 18624
rect 560294 18612 560300 18624
rect 174044 18584 560300 18612
rect 174044 18572 174050 18584
rect 560294 18572 560300 18584
rect 560352 18572 560358 18624
rect 443730 17892 443736 17944
rect 443788 17932 443794 17944
rect 449158 17932 449164 17944
rect 443788 17904 449164 17932
rect 443788 17892 443794 17904
rect 449158 17892 449164 17904
rect 449216 17892 449222 17944
rect 288342 17688 288348 17740
rect 288400 17728 288406 17740
rect 297358 17728 297364 17740
rect 288400 17700 297364 17728
rect 288400 17688 288406 17700
rect 297358 17688 297364 17700
rect 297416 17688 297422 17740
rect 148226 17620 148232 17672
rect 148284 17660 148290 17672
rect 226334 17660 226340 17672
rect 148284 17632 226340 17660
rect 148284 17620 148290 17632
rect 226334 17620 226340 17632
rect 226392 17620 226398 17672
rect 294138 17620 294144 17672
rect 294196 17660 294202 17672
rect 312630 17660 312636 17672
rect 294196 17632 312636 17660
rect 294196 17620 294202 17632
rect 312630 17620 312636 17632
rect 312688 17620 312694 17672
rect 355594 17620 355600 17672
rect 355652 17660 355658 17672
rect 365714 17660 365720 17672
rect 355652 17632 365720 17660
rect 355652 17620 355658 17632
rect 365714 17620 365720 17632
rect 365772 17620 365778 17672
rect 367738 17620 367744 17672
rect 367796 17660 367802 17672
rect 377398 17660 377404 17672
rect 367796 17632 377404 17660
rect 367796 17620 367802 17632
rect 377398 17620 377404 17632
rect 377456 17620 377462 17672
rect 161842 17552 161848 17604
rect 161900 17592 161906 17604
rect 398926 17592 398932 17604
rect 161900 17564 398932 17592
rect 161900 17552 161906 17564
rect 398926 17552 398932 17564
rect 398984 17552 398990 17604
rect 164418 17484 164424 17536
rect 164476 17524 164482 17536
rect 436094 17524 436100 17536
rect 164476 17496 436100 17524
rect 164476 17484 164482 17496
rect 436094 17484 436100 17496
rect 436152 17484 436158 17536
rect 164326 17416 164332 17468
rect 164384 17456 164390 17468
rect 441614 17456 441620 17468
rect 164384 17428 441620 17456
rect 164384 17416 164390 17428
rect 441614 17416 441620 17428
rect 441672 17416 441678 17468
rect 165890 17348 165896 17400
rect 165948 17388 165954 17400
rect 462314 17388 462320 17400
rect 165948 17360 462320 17388
rect 165948 17348 165954 17360
rect 462314 17348 462320 17360
rect 462372 17348 462378 17400
rect 171318 17280 171324 17332
rect 171376 17320 171382 17332
rect 523034 17320 523040 17332
rect 171376 17292 523040 17320
rect 171376 17280 171382 17292
rect 523034 17280 523040 17292
rect 523092 17280 523098 17332
rect 171226 17212 171232 17264
rect 171284 17252 171290 17264
rect 527174 17252 527180 17264
rect 171284 17224 527180 17252
rect 171284 17212 171290 17224
rect 527174 17212 527180 17224
rect 527232 17212 527238 17264
rect 342254 16804 342260 16856
rect 342312 16844 342318 16856
rect 346394 16844 346400 16856
rect 342312 16816 346400 16844
rect 342312 16804 342318 16816
rect 346394 16804 346400 16816
rect 346452 16804 346458 16856
rect 304442 16260 304448 16312
rect 304500 16300 304506 16312
rect 308398 16300 308404 16312
rect 304500 16272 308404 16300
rect 304500 16260 304506 16272
rect 308398 16260 308404 16272
rect 308456 16260 308462 16312
rect 149606 15920 149612 15972
rect 149664 15960 149670 15972
rect 248414 15960 248420 15972
rect 149664 15932 248420 15960
rect 149664 15920 149670 15932
rect 248414 15920 248420 15932
rect 248472 15920 248478 15972
rect 323578 15920 323584 15972
rect 323636 15960 323642 15972
rect 333238 15960 333244 15972
rect 323636 15932 333244 15960
rect 323636 15920 323642 15932
rect 333238 15920 333244 15932
rect 333296 15920 333302 15972
rect 334802 15920 334808 15972
rect 334860 15960 334866 15972
rect 339034 15960 339040 15972
rect 334860 15932 339040 15960
rect 334860 15920 334866 15932
rect 339034 15920 339040 15932
rect 339092 15920 339098 15972
rect 342898 15920 342904 15972
rect 342956 15960 342962 15972
rect 347866 15960 347872 15972
rect 342956 15932 347872 15960
rect 342956 15920 342962 15932
rect 347866 15920 347872 15932
rect 347924 15920 347930 15972
rect 35986 15852 35992 15904
rect 36044 15892 36050 15904
rect 124858 15892 124864 15904
rect 36044 15864 124864 15892
rect 36044 15852 36050 15864
rect 124858 15852 124864 15864
rect 124916 15852 124922 15904
rect 176286 15852 176292 15904
rect 176344 15892 176350 15904
rect 411898 15892 411904 15904
rect 176344 15864 411904 15892
rect 176344 15852 176350 15864
rect 411898 15852 411904 15864
rect 411956 15852 411962 15904
rect 349798 15716 349804 15768
rect 349856 15756 349862 15768
rect 352282 15756 352288 15768
rect 349856 15728 352288 15756
rect 349856 15716 349862 15728
rect 352282 15716 352288 15728
rect 352340 15716 352346 15768
rect 452746 15580 452752 15632
rect 452804 15620 452810 15632
rect 458174 15620 458180 15632
rect 452804 15592 458180 15620
rect 452804 15580 452810 15592
rect 458174 15580 458180 15592
rect 458232 15580 458238 15632
rect 152090 15104 152096 15156
rect 152148 15144 152154 15156
rect 276106 15144 276112 15156
rect 152148 15116 276112 15144
rect 152148 15104 152154 15116
rect 276106 15104 276112 15116
rect 276164 15104 276170 15156
rect 152182 15036 152188 15088
rect 152240 15076 152246 15088
rect 279050 15076 279056 15088
rect 152240 15048 279056 15076
rect 152240 15036 152246 15048
rect 279050 15036 279056 15048
rect 279108 15036 279114 15088
rect 308490 15036 308496 15088
rect 308548 15076 308554 15088
rect 319806 15076 319812 15088
rect 308548 15048 319812 15076
rect 308548 15036 308554 15048
rect 319806 15036 319812 15048
rect 319864 15036 319870 15088
rect 339310 15036 339316 15088
rect 339368 15076 339374 15088
rect 342806 15076 342812 15088
rect 339368 15048 342812 15076
rect 339368 15036 339374 15048
rect 342806 15036 342812 15048
rect 342864 15036 342870 15088
rect 151998 14968 152004 15020
rect 152056 15008 152062 15020
rect 283098 15008 283104 15020
rect 152056 14980 283104 15008
rect 152056 14968 152062 14980
rect 283098 14968 283104 14980
rect 283156 14968 283162 15020
rect 300118 14968 300124 15020
rect 300176 15008 300182 15020
rect 314746 15008 314752 15020
rect 300176 14980 314752 15008
rect 300176 14968 300182 14980
rect 314746 14968 314752 14980
rect 314804 14968 314810 15020
rect 334618 14968 334624 15020
rect 334676 15008 334682 15020
rect 340230 15008 340236 15020
rect 334676 14980 340236 15008
rect 334676 14968 334682 14980
rect 340230 14968 340236 14980
rect 340288 14968 340294 15020
rect 365070 14968 365076 15020
rect 365128 15008 365134 15020
rect 370498 15008 370504 15020
rect 365128 14980 370504 15008
rect 365128 14968 365134 14980
rect 370498 14968 370504 14980
rect 370556 14968 370562 15020
rect 153562 14900 153568 14952
rect 153620 14940 153626 14952
rect 297266 14940 297272 14952
rect 153620 14912 297272 14940
rect 153620 14900 153626 14912
rect 297266 14900 297272 14912
rect 297324 14900 297330 14952
rect 304258 14900 304264 14952
rect 304316 14940 304322 14952
rect 320726 14940 320732 14952
rect 304316 14912 320732 14940
rect 304316 14900 304322 14912
rect 320726 14900 320732 14912
rect 320784 14900 320790 14952
rect 324958 14900 324964 14952
rect 325016 14940 325022 14952
rect 347130 14940 347136 14952
rect 325016 14912 347136 14940
rect 325016 14900 325022 14912
rect 347130 14900 347136 14912
rect 347188 14900 347194 14952
rect 160094 14832 160100 14884
rect 160152 14872 160158 14884
rect 384298 14872 384304 14884
rect 160152 14844 384304 14872
rect 160152 14832 160158 14844
rect 384298 14832 384304 14844
rect 384356 14832 384362 14884
rect 160186 14764 160192 14816
rect 160244 14804 160250 14816
rect 387794 14804 387800 14816
rect 160244 14776 387800 14804
rect 160244 14764 160250 14776
rect 387794 14764 387800 14776
rect 387852 14764 387858 14816
rect 160278 14696 160284 14748
rect 160336 14736 160342 14748
rect 390646 14736 390652 14748
rect 160336 14708 390652 14736
rect 160336 14696 160342 14708
rect 390646 14696 390652 14708
rect 390704 14696 390710 14748
rect 161750 14628 161756 14680
rect 161808 14668 161814 14680
rect 400858 14668 400864 14680
rect 161808 14640 400864 14668
rect 161808 14628 161814 14640
rect 400858 14628 400864 14640
rect 400916 14628 400922 14680
rect 162854 14560 162860 14612
rect 162912 14600 162918 14612
rect 420914 14600 420920 14612
rect 162912 14572 420920 14600
rect 162912 14560 162918 14572
rect 420914 14560 420920 14572
rect 420972 14560 420978 14612
rect 449158 14560 449164 14612
rect 449216 14600 449222 14612
rect 454586 14600 454592 14612
rect 449216 14572 454592 14600
rect 449216 14560 449222 14572
rect 454586 14560 454592 14572
rect 454644 14560 454650 14612
rect 165798 14492 165804 14544
rect 165856 14532 165862 14544
rect 459186 14532 459192 14544
rect 165856 14504 459192 14532
rect 165856 14492 165862 14504
rect 459186 14492 459192 14504
rect 459244 14492 459250 14544
rect 468478 14492 468484 14544
rect 468536 14532 468542 14544
rect 482278 14532 482284 14544
rect 468536 14504 482284 14532
rect 468536 14492 468542 14504
rect 482278 14492 482284 14504
rect 482336 14492 482342 14544
rect 174814 14424 174820 14476
rect 174872 14464 174878 14476
rect 567562 14464 567568 14476
rect 174872 14436 567568 14464
rect 174872 14424 174878 14436
rect 567562 14424 567568 14436
rect 567620 14424 567626 14476
rect 150802 14356 150808 14408
rect 150860 14396 150866 14408
rect 264974 14396 264980 14408
rect 150860 14368 264980 14396
rect 150860 14356 150866 14368
rect 264974 14356 264980 14368
rect 265032 14356 265038 14408
rect 348418 14356 348424 14408
rect 348476 14396 348482 14408
rect 350902 14396 350908 14408
rect 348476 14368 350908 14396
rect 348476 14356 348482 14368
rect 350902 14356 350908 14368
rect 350960 14356 350966 14408
rect 150710 14288 150716 14340
rect 150768 14328 150774 14340
rect 261754 14328 261760 14340
rect 150768 14300 261760 14328
rect 150768 14288 150774 14300
rect 261754 14288 261760 14300
rect 261812 14288 261818 14340
rect 147030 14220 147036 14272
rect 147088 14260 147094 14272
rect 190454 14260 190460 14272
rect 147088 14232 190460 14260
rect 147088 14220 147094 14232
rect 190454 14220 190460 14232
rect 190512 14220 190518 14272
rect 364978 13880 364984 13932
rect 365036 13920 365042 13932
rect 367738 13920 367744 13932
rect 365036 13892 367744 13920
rect 365036 13880 365042 13892
rect 367738 13880 367744 13892
rect 367796 13880 367802 13932
rect 319438 13812 319444 13864
rect 319496 13852 319502 13864
rect 322198 13852 322204 13864
rect 319496 13824 322204 13852
rect 319496 13812 319502 13824
rect 322198 13812 322204 13824
rect 322256 13812 322262 13864
rect 321186 13744 321192 13796
rect 321244 13784 321250 13796
rect 326338 13784 326344 13796
rect 321244 13756 326344 13784
rect 321244 13744 321250 13756
rect 326338 13744 326344 13756
rect 326396 13744 326402 13796
rect 353938 13744 353944 13796
rect 353996 13784 354002 13796
rect 356698 13784 356704 13796
rect 353996 13756 356704 13784
rect 353996 13744 354002 13756
rect 356698 13744 356704 13756
rect 356756 13744 356762 13796
rect 479518 13744 479524 13796
rect 479576 13784 479582 13796
rect 481726 13784 481732 13796
rect 479576 13756 481732 13784
rect 479576 13744 479582 13756
rect 481726 13744 481732 13756
rect 481784 13744 481790 13796
rect 341518 13676 341524 13728
rect 341576 13716 341582 13728
rect 347038 13716 347044 13728
rect 341576 13688 347044 13716
rect 341576 13676 341582 13688
rect 347038 13676 347044 13688
rect 347096 13676 347102 13728
rect 329098 13200 329104 13252
rect 329156 13240 329162 13252
rect 334618 13240 334624 13252
rect 329156 13212 334624 13240
rect 329156 13200 329162 13212
rect 334618 13200 334624 13212
rect 334676 13200 334682 13252
rect 493318 13064 493324 13116
rect 493376 13104 493382 13116
rect 507854 13104 507860 13116
rect 493376 13076 507860 13104
rect 493376 13064 493382 13076
rect 507854 13064 507860 13076
rect 507912 13064 507918 13116
rect 340046 12452 340052 12504
rect 340104 12492 340110 12504
rect 342990 12492 342996 12504
rect 340104 12464 342996 12492
rect 340104 12452 340110 12464
rect 342990 12452 342996 12464
rect 343048 12452 343054 12504
rect 146386 12384 146392 12436
rect 146444 12424 146450 12436
rect 214466 12424 214472 12436
rect 146444 12396 214472 12424
rect 146444 12384 146450 12396
rect 214466 12384 214472 12396
rect 214524 12384 214530 12436
rect 358078 12384 358084 12436
rect 358136 12424 358142 12436
rect 361574 12424 361580 12436
rect 358136 12396 361580 12424
rect 358136 12384 358142 12396
rect 361574 12384 361580 12396
rect 361632 12384 361638 12436
rect 458818 12384 458824 12436
rect 458876 12424 458882 12436
rect 461670 12424 461676 12436
rect 458876 12396 461676 12424
rect 458876 12384 458882 12396
rect 461670 12384 461676 12396
rect 461728 12384 461734 12436
rect 148134 12316 148140 12368
rect 148192 12356 148198 12368
rect 222746 12356 222752 12368
rect 148192 12328 222752 12356
rect 148192 12316 148198 12328
rect 222746 12316 222752 12328
rect 222804 12316 222810 12368
rect 147950 12248 147956 12300
rect 148008 12288 148014 12300
rect 226426 12288 226432 12300
rect 148008 12260 226432 12288
rect 148008 12248 148014 12260
rect 226426 12248 226432 12260
rect 226484 12248 226490 12300
rect 307110 12248 307116 12300
rect 307168 12288 307174 12300
rect 311894 12288 311900 12300
rect 307168 12260 311900 12288
rect 307168 12248 307174 12260
rect 311894 12248 311900 12260
rect 311952 12248 311958 12300
rect 148042 12180 148048 12232
rect 148100 12220 148106 12232
rect 229370 12220 229376 12232
rect 148100 12192 229376 12220
rect 148100 12180 148106 12192
rect 229370 12180 229376 12192
rect 229428 12180 229434 12232
rect 149514 12112 149520 12164
rect 149572 12152 149578 12164
rect 240134 12152 240140 12164
rect 149572 12124 240140 12152
rect 149572 12112 149578 12124
rect 240134 12112 240140 12124
rect 240192 12112 240198 12164
rect 320726 12112 320732 12164
rect 320784 12152 320790 12164
rect 320784 12124 325694 12152
rect 320784 12112 320790 12124
rect 149422 12044 149428 12096
rect 149480 12084 149486 12096
rect 242894 12084 242900 12096
rect 149480 12056 242900 12084
rect 149480 12044 149486 12056
rect 242894 12044 242900 12056
rect 242952 12044 242958 12096
rect 319622 12044 319628 12096
rect 319680 12084 319686 12096
rect 322290 12084 322296 12096
rect 319680 12056 322296 12084
rect 319680 12044 319686 12056
rect 322290 12044 322296 12056
rect 322348 12044 322354 12096
rect 325666 12084 325694 12124
rect 352650 12112 352656 12164
rect 352708 12152 352714 12164
rect 357526 12152 357532 12164
rect 352708 12124 357532 12152
rect 352708 12112 352714 12124
rect 357526 12112 357532 12124
rect 357584 12112 357590 12164
rect 329098 12084 329104 12096
rect 325666 12056 329104 12084
rect 329098 12044 329104 12056
rect 329156 12044 329162 12096
rect 347866 12044 347872 12096
rect 347924 12084 347930 12096
rect 359458 12084 359464 12096
rect 347924 12056 359464 12084
rect 347924 12044 347930 12056
rect 359458 12044 359464 12056
rect 359516 12044 359522 12096
rect 165154 11976 165160 12028
rect 165212 12016 165218 12028
rect 382366 12016 382372 12028
rect 165212 11988 382372 12016
rect 165212 11976 165218 11988
rect 382366 11976 382372 11988
rect 382424 11976 382430 12028
rect 382918 11976 382924 12028
rect 382976 12016 382982 12028
rect 389818 12016 389824 12028
rect 382976 11988 389824 12016
rect 382976 11976 382982 11988
rect 389818 11976 389824 11988
rect 389876 11976 389882 12028
rect 161658 11908 161664 11960
rect 161716 11948 161722 11960
rect 402514 11948 402520 11960
rect 161716 11920 402520 11948
rect 161716 11908 161722 11920
rect 402514 11908 402520 11920
rect 402572 11908 402578 11960
rect 161566 11840 161572 11892
rect 161624 11880 161630 11892
rect 406010 11880 406016 11892
rect 161624 11852 406016 11880
rect 161624 11840 161630 11852
rect 406010 11840 406016 11852
rect 406068 11840 406074 11892
rect 165706 11772 165712 11824
rect 165764 11812 165770 11824
rect 455690 11812 455696 11824
rect 165764 11784 455696 11812
rect 165764 11772 165770 11784
rect 455690 11772 455696 11784
rect 455748 11772 455754 11824
rect 476758 11772 476764 11824
rect 476816 11812 476822 11824
rect 479518 11812 479524 11824
rect 476816 11784 479524 11812
rect 476816 11772 476822 11784
rect 479518 11772 479524 11784
rect 479576 11772 479582 11824
rect 126974 11704 126980 11756
rect 127032 11744 127038 11756
rect 128170 11744 128176 11756
rect 127032 11716 128176 11744
rect 127032 11704 127038 11716
rect 128170 11704 128176 11716
rect 128228 11704 128234 11756
rect 135254 11704 135260 11756
rect 135312 11744 135318 11756
rect 136450 11744 136456 11756
rect 135312 11716 136456 11744
rect 135312 11704 135318 11716
rect 136450 11704 136456 11716
rect 136508 11704 136514 11756
rect 169846 11704 169852 11756
rect 169904 11744 169910 11756
rect 511258 11744 511264 11756
rect 169904 11716 511264 11744
rect 169904 11704 169910 11716
rect 511258 11704 511264 11716
rect 511316 11704 511322 11756
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 226334 11636 226340 11688
rect 226392 11676 226398 11688
rect 227530 11676 227536 11688
rect 226392 11648 227536 11676
rect 226392 11636 226398 11648
rect 227530 11636 227536 11648
rect 227588 11636 227594 11688
rect 259454 11636 259460 11688
rect 259512 11676 259518 11688
rect 260650 11676 260656 11688
rect 259512 11648 260656 11676
rect 259512 11636 259518 11648
rect 260650 11636 260656 11648
rect 260708 11636 260714 11688
rect 311158 11636 311164 11688
rect 311216 11676 311222 11688
rect 314654 11676 314660 11688
rect 311216 11648 314660 11676
rect 311216 11636 311222 11648
rect 314654 11636 314660 11648
rect 314712 11636 314718 11688
rect 327718 11636 327724 11688
rect 327776 11676 327782 11688
rect 330478 11676 330484 11688
rect 327776 11648 330484 11676
rect 327776 11636 327782 11648
rect 330478 11636 330484 11648
rect 330536 11636 330542 11688
rect 316678 10956 316684 11008
rect 316736 10996 316742 11008
rect 319438 10996 319444 11008
rect 316736 10968 319444 10996
rect 316736 10956 316742 10968
rect 319438 10956 319444 10968
rect 319496 10956 319502 11008
rect 339034 10956 339040 11008
rect 339092 10996 339098 11008
rect 342714 10996 342720 11008
rect 339092 10968 342720 10996
rect 339092 10956 339098 10968
rect 342714 10956 342720 10968
rect 342772 10956 342778 11008
rect 347130 10956 347136 11008
rect 347188 10996 347194 11008
rect 349246 10996 349252 11008
rect 347188 10968 349252 10996
rect 347188 10956 347194 10968
rect 349246 10956 349252 10968
rect 349304 10956 349310 11008
rect 318058 10888 318064 10940
rect 318116 10928 318122 10940
rect 322382 10928 322388 10940
rect 318116 10900 322388 10928
rect 318116 10888 318122 10900
rect 322382 10888 322388 10900
rect 322440 10888 322446 10940
rect 112346 10684 112352 10736
rect 112404 10724 112410 10736
rect 138382 10724 138388 10736
rect 112404 10696 138388 10724
rect 112404 10684 112410 10696
rect 138382 10684 138388 10696
rect 138440 10684 138446 10736
rect 92474 10616 92480 10668
rect 92532 10656 92538 10668
rect 130378 10656 130384 10668
rect 92532 10628 130384 10656
rect 92532 10616 92538 10628
rect 130378 10616 130384 10628
rect 130436 10616 130442 10668
rect 89162 10548 89168 10600
rect 89220 10588 89226 10600
rect 137002 10588 137008 10600
rect 89220 10560 137008 10588
rect 89220 10548 89226 10560
rect 137002 10548 137008 10560
rect 137060 10548 137066 10600
rect 74994 10480 75000 10532
rect 75052 10520 75058 10532
rect 134518 10520 134524 10532
rect 75052 10492 134524 10520
rect 75052 10480 75058 10492
rect 134518 10480 134524 10492
rect 134576 10480 134582 10532
rect 71498 10412 71504 10464
rect 71556 10452 71562 10464
rect 135898 10452 135904 10464
rect 71556 10424 135904 10452
rect 71556 10412 71562 10424
rect 135898 10412 135904 10424
rect 135956 10412 135962 10464
rect 20162 10344 20168 10396
rect 20220 10384 20226 10396
rect 95878 10384 95884 10396
rect 20220 10356 95884 10384
rect 20220 10344 20226 10356
rect 95878 10344 95884 10356
rect 95936 10344 95942 10396
rect 106458 10344 106464 10396
rect 106516 10384 106522 10396
rect 138474 10384 138480 10396
rect 106516 10356 138480 10384
rect 106516 10344 106522 10356
rect 138474 10344 138480 10356
rect 138532 10344 138538 10396
rect 350902 10344 350908 10396
rect 350960 10384 350966 10396
rect 363506 10384 363512 10396
rect 350960 10356 363512 10384
rect 350960 10344 350966 10356
rect 363506 10344 363512 10356
rect 363564 10344 363570 10396
rect 365714 10344 365720 10396
rect 365772 10384 365778 10396
rect 374086 10384 374092 10396
rect 365772 10356 374092 10384
rect 365772 10344 365778 10356
rect 374086 10344 374092 10356
rect 374144 10344 374150 10396
rect 458174 10344 458180 10396
rect 458232 10384 458238 10396
rect 465718 10384 465724 10396
rect 458232 10356 465724 10384
rect 458232 10344 458238 10356
rect 465718 10344 465724 10356
rect 465776 10344 465782 10396
rect 56778 10276 56784 10328
rect 56836 10316 56842 10328
rect 134334 10316 134340 10328
rect 56836 10288 134340 10316
rect 56836 10276 56842 10288
rect 134334 10276 134340 10288
rect 134392 10276 134398 10328
rect 169754 10276 169760 10328
rect 169812 10316 169818 10328
rect 503714 10316 503720 10328
rect 169812 10288 503720 10316
rect 169812 10276 169818 10288
rect 503714 10276 503720 10288
rect 503772 10276 503778 10328
rect 307202 9596 307208 9648
rect 307260 9636 307266 9648
rect 309318 9636 309324 9648
rect 307260 9608 309324 9636
rect 307260 9596 307266 9608
rect 309318 9596 309324 9608
rect 309376 9596 309382 9648
rect 320910 9596 320916 9648
rect 320968 9636 320974 9648
rect 324682 9636 324688 9648
rect 320968 9608 324688 9636
rect 320968 9596 320974 9608
rect 324682 9596 324688 9608
rect 324740 9596 324746 9648
rect 335998 9596 336004 9648
rect 336056 9636 336062 9648
rect 342162 9636 342168 9648
rect 336056 9608 342168 9636
rect 336056 9596 336062 9608
rect 342162 9596 342168 9608
rect 342220 9596 342226 9648
rect 320818 9528 320824 9580
rect 320876 9568 320882 9580
rect 324774 9568 324780 9580
rect 320876 9540 324780 9568
rect 320876 9528 320882 9540
rect 324774 9528 324780 9540
rect 324832 9528 324838 9580
rect 109310 9392 109316 9444
rect 109368 9432 109374 9444
rect 138290 9432 138296 9444
rect 109368 9404 138296 9432
rect 109368 9392 109374 9404
rect 138290 9392 138296 9404
rect 138348 9392 138354 9444
rect 82078 9324 82084 9376
rect 82136 9364 82142 9376
rect 136910 9364 136916 9376
rect 82136 9336 136916 9364
rect 82136 9324 82142 9336
rect 136910 9324 136916 9336
rect 136968 9324 136974 9376
rect 77386 9256 77392 9308
rect 77444 9296 77450 9308
rect 135714 9296 135720 9308
rect 77444 9268 135720 9296
rect 77444 9256 77450 9268
rect 135714 9256 135720 9268
rect 135772 9256 135778 9308
rect 73798 9188 73804 9240
rect 73856 9228 73862 9240
rect 135622 9228 135628 9240
rect 73856 9200 135628 9228
rect 73856 9188 73862 9200
rect 135622 9188 135628 9200
rect 135680 9188 135686 9240
rect 177482 9188 177488 9240
rect 177540 9228 177546 9240
rect 207382 9228 207388 9240
rect 177540 9200 207388 9228
rect 177540 9188 177546 9200
rect 207382 9188 207388 9200
rect 207440 9188 207446 9240
rect 70302 9120 70308 9172
rect 70360 9160 70366 9172
rect 135806 9160 135812 9172
rect 70360 9132 135812 9160
rect 70360 9120 70366 9132
rect 135806 9120 135812 9132
rect 135864 9120 135870 9172
rect 146294 9120 146300 9172
rect 146352 9160 146358 9172
rect 210970 9160 210976 9172
rect 146352 9132 210976 9160
rect 146352 9120 146358 9132
rect 210970 9120 210976 9132
rect 211028 9120 211034 9172
rect 352282 9120 352288 9172
rect 352340 9160 352346 9172
rect 364610 9160 364616 9172
rect 352340 9132 364616 9160
rect 352340 9120 352346 9132
rect 364610 9120 364616 9132
rect 364668 9120 364674 9172
rect 43070 9052 43076 9104
rect 43128 9092 43134 9104
rect 122098 9092 122104 9104
rect 43128 9064 122104 9092
rect 43128 9052 43134 9064
rect 122098 9052 122104 9064
rect 122156 9052 122162 9104
rect 149330 9052 149336 9104
rect 149388 9092 149394 9104
rect 247586 9092 247592 9104
rect 149388 9064 247592 9092
rect 149388 9052 149394 9064
rect 247586 9052 247592 9064
rect 247644 9052 247650 9104
rect 282178 9052 282184 9104
rect 282236 9092 282242 9104
rect 302142 9092 302148 9104
rect 282236 9064 302148 9092
rect 282236 9052 282242 9064
rect 302142 9052 302148 9064
rect 302200 9052 302206 9104
rect 304350 9052 304356 9104
rect 304408 9092 304414 9104
rect 312262 9092 312268 9104
rect 304408 9064 312268 9092
rect 304408 9052 304414 9064
rect 312262 9052 312268 9064
rect 312320 9052 312326 9104
rect 315298 9052 315304 9104
rect 315356 9092 315362 9104
rect 330754 9092 330760 9104
rect 315356 9064 330760 9092
rect 315356 9052 315362 9064
rect 330754 9052 330760 9064
rect 330812 9052 330818 9104
rect 338758 9052 338764 9104
rect 338816 9092 338822 9104
rect 351454 9092 351460 9104
rect 338816 9064 351460 9092
rect 338816 9052 338822 9064
rect 351454 9052 351460 9064
rect 351512 9052 351518 9104
rect 361574 9052 361580 9104
rect 361632 9092 361638 9104
rect 377674 9092 377680 9104
rect 361632 9064 377680 9092
rect 361632 9052 361638 9064
rect 377674 9052 377680 9064
rect 377732 9052 377738 9104
rect 53742 8984 53748 9036
rect 53800 9024 53806 9036
rect 134242 9024 134248 9036
rect 53800 8996 134248 9024
rect 53800 8984 53806 8996
rect 134242 8984 134248 8996
rect 134300 8984 134306 9036
rect 161474 8984 161480 9036
rect 161532 9024 161538 9036
rect 407206 9024 407212 9036
rect 161532 8996 407212 9024
rect 161532 8984 161538 8996
rect 407206 8984 407212 8996
rect 407264 8984 407270 9036
rect 14734 8916 14740 8968
rect 14792 8956 14798 8968
rect 131758 8956 131764 8968
rect 14792 8928 131764 8956
rect 14792 8916 14798 8928
rect 131758 8916 131764 8928
rect 131816 8916 131822 8968
rect 168466 8916 168472 8968
rect 168524 8956 168530 8968
rect 493502 8956 493508 8968
rect 168524 8928 493508 8956
rect 168524 8916 168530 8928
rect 493502 8916 493508 8928
rect 493560 8916 493566 8968
rect 507854 8916 507860 8968
rect 507912 8956 507918 8968
rect 526622 8956 526628 8968
rect 507912 8928 526628 8956
rect 507912 8916 507918 8928
rect 526622 8916 526628 8928
rect 526680 8916 526686 8968
rect 312630 8304 312636 8356
rect 312688 8344 312694 8356
rect 316218 8344 316224 8356
rect 312688 8316 316224 8344
rect 312688 8304 312694 8316
rect 316218 8304 316224 8316
rect 316276 8304 316282 8356
rect 297358 8236 297364 8288
rect 297416 8276 297422 8288
rect 303522 8276 303528 8288
rect 297416 8248 303528 8276
rect 297416 8236 297422 8248
rect 303522 8236 303528 8248
rect 303580 8236 303586 8288
rect 377398 8236 377404 8288
rect 377456 8276 377462 8288
rect 379974 8276 379980 8288
rect 377456 8248 379980 8276
rect 377456 8236 377462 8248
rect 379974 8236 379980 8248
rect 380032 8236 380038 8288
rect 135254 8100 135260 8152
rect 135312 8140 135318 8152
rect 135438 8140 135444 8152
rect 135312 8112 135444 8140
rect 135312 8100 135318 8112
rect 135438 8100 135444 8112
rect 135496 8100 135502 8152
rect 123478 7896 123484 7948
rect 123536 7936 123542 7948
rect 139578 7936 139584 7948
rect 123536 7908 139584 7936
rect 123536 7896 123542 7908
rect 139578 7896 139584 7908
rect 139636 7896 139642 7948
rect 66714 7828 66720 7880
rect 66772 7868 66778 7880
rect 135530 7868 135536 7880
rect 66772 7840 135536 7868
rect 66772 7828 66778 7840
rect 135530 7828 135536 7840
rect 135588 7828 135594 7880
rect 52546 7760 52552 7812
rect 52604 7800 52610 7812
rect 134058 7800 134064 7812
rect 52604 7772 134064 7800
rect 52604 7760 52610 7772
rect 134058 7760 134064 7772
rect 134116 7760 134122 7812
rect 50154 7692 50160 7744
rect 50212 7732 50218 7744
rect 134150 7732 134156 7744
rect 50212 7704 134156 7732
rect 50212 7692 50218 7704
rect 134150 7692 134156 7704
rect 134208 7692 134214 7744
rect 312538 7692 312544 7744
rect 312596 7732 312602 7744
rect 323302 7732 323308 7744
rect 312596 7704 323308 7732
rect 312596 7692 312602 7704
rect 323302 7692 323308 7704
rect 323360 7692 323366 7744
rect 28902 7624 28908 7676
rect 28960 7664 28966 7676
rect 126330 7664 126336 7676
rect 28960 7636 126336 7664
rect 28960 7624 28966 7636
rect 126330 7624 126336 7636
rect 126388 7624 126394 7676
rect 314746 7624 314752 7676
rect 314804 7664 314810 7676
rect 327074 7664 327080 7676
rect 314804 7636 327080 7664
rect 314804 7624 314810 7636
rect 327074 7624 327080 7636
rect 327132 7624 327138 7676
rect 334710 7624 334716 7676
rect 334768 7664 334774 7676
rect 356330 7664 356336 7676
rect 334768 7636 356336 7664
rect 334768 7624 334774 7636
rect 356330 7624 356336 7636
rect 356388 7624 356394 7676
rect 15930 7556 15936 7608
rect 15988 7596 15994 7608
rect 131666 7596 131672 7608
rect 15988 7568 131672 7596
rect 15988 7556 15994 7568
rect 131666 7556 131672 7568
rect 131724 7556 131730 7608
rect 164234 7556 164240 7608
rect 164292 7596 164298 7608
rect 443822 7596 443828 7608
rect 164292 7568 443828 7596
rect 164292 7556 164298 7568
rect 443822 7556 443828 7568
rect 443880 7556 443886 7608
rect 454586 7556 454592 7608
rect 454644 7596 454650 7608
rect 473446 7596 473452 7608
rect 454644 7568 473452 7596
rect 454644 7556 454650 7568
rect 473446 7556 473452 7568
rect 473504 7556 473510 7608
rect 311894 7488 311900 7540
rect 311952 7528 311958 7540
rect 317414 7528 317420 7540
rect 311952 7500 317420 7528
rect 311952 7488 311958 7500
rect 317414 7488 317420 7500
rect 317472 7488 317478 7540
rect 149974 6808 149980 6860
rect 150032 6848 150038 6860
rect 203886 6848 203892 6860
rect 150032 6820 203892 6848
rect 150032 6808 150038 6820
rect 203886 6808 203892 6820
rect 203944 6808 203950 6860
rect 149238 6740 149244 6792
rect 149296 6780 149302 6792
rect 246390 6780 246396 6792
rect 149296 6752 246396 6780
rect 149296 6740 149302 6752
rect 246390 6740 246396 6752
rect 246448 6740 246454 6792
rect 150618 6672 150624 6724
rect 150676 6712 150682 6724
rect 267734 6712 267740 6724
rect 150676 6684 267740 6712
rect 150676 6672 150682 6684
rect 267734 6672 267740 6684
rect 267792 6672 267798 6724
rect 151814 6604 151820 6656
rect 151872 6644 151878 6656
rect 278314 6644 278320 6656
rect 151872 6616 278320 6644
rect 151872 6604 151878 6616
rect 278314 6604 278320 6616
rect 278372 6604 278378 6656
rect 40678 6536 40684 6588
rect 40736 6576 40742 6588
rect 132678 6576 132684 6588
rect 40736 6548 132684 6576
rect 40736 6536 40742 6548
rect 132678 6536 132684 6548
rect 132736 6536 132742 6588
rect 151906 6536 151912 6588
rect 151964 6576 151970 6588
rect 281902 6576 281908 6588
rect 151964 6548 281908 6576
rect 151964 6536 151970 6548
rect 281902 6536 281908 6548
rect 281960 6536 281966 6588
rect 333238 6536 333244 6588
rect 333296 6576 333302 6588
rect 338666 6576 338672 6588
rect 333296 6548 338672 6576
rect 333296 6536 333302 6548
rect 338666 6536 338672 6548
rect 338724 6536 338730 6588
rect 38378 6468 38384 6520
rect 38436 6508 38442 6520
rect 133046 6508 133052 6520
rect 38436 6480 133052 6508
rect 38436 6468 38442 6480
rect 133046 6468 133052 6480
rect 133104 6468 133110 6520
rect 153470 6468 153476 6520
rect 153528 6508 153534 6520
rect 292574 6508 292580 6520
rect 153528 6480 292580 6508
rect 153528 6468 153534 6480
rect 292574 6468 292580 6480
rect 292632 6468 292638 6520
rect 324682 6468 324688 6520
rect 324740 6508 324746 6520
rect 334066 6508 334072 6520
rect 324740 6480 334072 6508
rect 324740 6468 324746 6480
rect 334066 6468 334072 6480
rect 334124 6468 334130 6520
rect 37182 6400 37188 6452
rect 37240 6440 37246 6452
rect 132770 6440 132776 6452
rect 37240 6412 132776 6440
rect 37240 6400 37246 6412
rect 132770 6400 132776 6412
rect 132828 6400 132834 6452
rect 153378 6400 153384 6452
rect 153436 6440 153442 6452
rect 296070 6440 296076 6452
rect 153436 6412 296076 6440
rect 153436 6400 153442 6412
rect 296070 6400 296076 6412
rect 296128 6400 296134 6452
rect 324774 6400 324780 6452
rect 324832 6440 324838 6452
rect 333974 6440 333980 6452
rect 324832 6412 333980 6440
rect 324832 6400 324838 6412
rect 333974 6400 333980 6412
rect 334032 6400 334038 6452
rect 340230 6400 340236 6452
rect 340288 6440 340294 6452
rect 352834 6440 352840 6452
rect 340288 6412 352840 6440
rect 340288 6400 340294 6412
rect 352834 6400 352840 6412
rect 352892 6400 352898 6452
rect 33594 6332 33600 6384
rect 33652 6372 33658 6384
rect 132954 6372 132960 6384
rect 33652 6344 132960 6372
rect 33652 6332 33658 6344
rect 132954 6332 132960 6344
rect 133012 6332 133018 6384
rect 153286 6332 153292 6384
rect 153344 6372 153350 6384
rect 299658 6372 299664 6384
rect 153344 6344 299664 6372
rect 153344 6332 153350 6344
rect 299658 6332 299664 6344
rect 299716 6332 299722 6384
rect 330754 6332 330760 6384
rect 330812 6372 330818 6384
rect 343634 6372 343640 6384
rect 330812 6344 343640 6372
rect 330812 6332 330818 6344
rect 343634 6332 343640 6344
rect 343692 6332 343698 6384
rect 31294 6264 31300 6316
rect 31352 6304 31358 6316
rect 133138 6304 133144 6316
rect 31352 6276 133144 6304
rect 31352 6264 31358 6276
rect 133138 6264 133144 6276
rect 133196 6264 133202 6316
rect 153194 6264 153200 6316
rect 153252 6304 153258 6316
rect 300762 6304 300768 6316
rect 153252 6276 300768 6304
rect 153252 6264 153258 6276
rect 300762 6264 300768 6276
rect 300820 6264 300826 6316
rect 305638 6264 305644 6316
rect 305696 6304 305702 6316
rect 309226 6304 309232 6316
rect 305696 6276 309232 6304
rect 305696 6264 305702 6276
rect 309226 6264 309232 6276
rect 309284 6264 309290 6316
rect 309318 6264 309324 6316
rect 309376 6304 309382 6316
rect 339862 6304 339868 6316
rect 309376 6276 339868 6304
rect 309376 6264 309382 6276
rect 339862 6264 339868 6276
rect 339920 6264 339926 6316
rect 342990 6264 342996 6316
rect 343048 6304 343054 6316
rect 357158 6304 357164 6316
rect 343048 6276 357164 6304
rect 343048 6264 343054 6276
rect 357158 6264 357164 6276
rect 357216 6264 357222 6316
rect 30098 6196 30104 6248
rect 30156 6236 30162 6248
rect 132862 6236 132868 6248
rect 30156 6208 132868 6236
rect 30156 6196 30162 6208
rect 132862 6196 132868 6208
rect 132920 6196 132926 6248
rect 175182 6196 175188 6248
rect 175240 6236 175246 6248
rect 573910 6236 573916 6248
rect 175240 6208 573916 6236
rect 175240 6196 175246 6208
rect 573910 6196 573916 6208
rect 573968 6196 573974 6248
rect 24210 6128 24216 6180
rect 24268 6168 24274 6180
rect 131574 6168 131580 6180
rect 24268 6140 131580 6168
rect 24268 6128 24274 6140
rect 131574 6128 131580 6140
rect 131632 6128 131638 6180
rect 176562 6128 176568 6180
rect 176620 6168 176626 6180
rect 578602 6168 578608 6180
rect 176620 6140 578608 6168
rect 176620 6128 176626 6140
rect 578602 6128 578608 6140
rect 578660 6128 578666 6180
rect 144914 6060 144920 6112
rect 144972 6100 144978 6112
rect 196802 6100 196808 6112
rect 144972 6072 196808 6100
rect 144972 6060 144978 6072
rect 196802 6060 196808 6072
rect 196860 6060 196866 6112
rect 356698 5924 356704 5976
rect 356756 5964 356762 5976
rect 362954 5964 362960 5976
rect 356756 5936 362960 5964
rect 356756 5924 356762 5936
rect 362954 5924 362960 5936
rect 363012 5924 363018 5976
rect 351454 5856 351460 5908
rect 351512 5896 351518 5908
rect 353294 5896 353300 5908
rect 351512 5868 353300 5896
rect 351512 5856 351518 5868
rect 353294 5856 353300 5868
rect 353352 5856 353358 5908
rect 319530 5516 319536 5568
rect 319588 5556 319594 5568
rect 324406 5556 324412 5568
rect 319588 5528 324412 5556
rect 319588 5516 319594 5528
rect 324406 5516 324412 5528
rect 324464 5516 324470 5568
rect 326338 5516 326344 5568
rect 326396 5556 326402 5568
rect 332686 5556 332692 5568
rect 326396 5528 332692 5556
rect 326396 5516 326402 5528
rect 332686 5516 332692 5528
rect 332744 5516 332750 5568
rect 479518 5516 479524 5568
rect 479576 5556 479582 5568
rect 482830 5556 482836 5568
rect 479576 5528 482836 5556
rect 479576 5516 479582 5528
rect 482830 5516 482836 5528
rect 482888 5516 482894 5568
rect 143810 5380 143816 5432
rect 143868 5420 143874 5432
rect 149238 5420 149244 5432
rect 143868 5392 149244 5420
rect 143868 5380 143874 5392
rect 149238 5380 149244 5392
rect 149296 5380 149302 5432
rect 122282 5312 122288 5364
rect 122340 5352 122346 5364
rect 139946 5352 139952 5364
rect 122340 5324 139952 5352
rect 122340 5312 122346 5324
rect 139946 5312 139952 5324
rect 140004 5312 140010 5364
rect 110506 5244 110512 5296
rect 110564 5284 110570 5296
rect 129182 5284 129188 5296
rect 110564 5256 129188 5284
rect 110564 5244 110570 5256
rect 129182 5244 129188 5256
rect 129240 5244 129246 5296
rect 108114 5176 108120 5228
rect 108172 5216 108178 5228
rect 138198 5216 138204 5228
rect 108172 5188 138204 5216
rect 108172 5176 108178 5188
rect 138198 5176 138204 5188
rect 138256 5176 138262 5228
rect 142338 5176 142344 5228
rect 142396 5216 142402 5228
rect 155402 5216 155408 5228
rect 142396 5188 155408 5216
rect 142396 5176 142402 5188
rect 155402 5176 155408 5188
rect 155460 5176 155466 5228
rect 104526 5108 104532 5160
rect 104584 5148 104590 5160
rect 138934 5148 138940 5160
rect 104584 5120 138940 5148
rect 104584 5108 104590 5120
rect 138934 5108 138940 5120
rect 138992 5108 138998 5160
rect 142430 5108 142436 5160
rect 142488 5148 142494 5160
rect 157794 5148 157800 5160
rect 142488 5120 157800 5148
rect 142488 5108 142494 5120
rect 157794 5108 157800 5120
rect 157852 5108 157858 5160
rect 56042 5040 56048 5092
rect 56100 5080 56106 5092
rect 134426 5080 134432 5092
rect 56100 5052 134432 5080
rect 56100 5040 56106 5052
rect 134426 5040 134432 5052
rect 134484 5040 134490 5092
rect 143902 5040 143908 5092
rect 143960 5080 143966 5092
rect 169570 5080 169576 5092
rect 143960 5052 169576 5080
rect 143960 5040 143966 5052
rect 169570 5040 169576 5052
rect 169628 5040 169634 5092
rect 23014 4972 23020 5024
rect 23072 5012 23078 5024
rect 131390 5012 131396 5024
rect 23072 4984 131396 5012
rect 23072 4972 23078 4984
rect 131390 4972 131396 4984
rect 131448 4972 131454 5024
rect 143994 4972 144000 5024
rect 144052 5012 144058 5024
rect 173158 5012 173164 5024
rect 144052 4984 173164 5012
rect 144052 4972 144058 4984
rect 173158 4972 173164 4984
rect 173216 4972 173222 5024
rect 220446 5012 220452 5024
rect 200086 4984 220452 5012
rect 19426 4904 19432 4956
rect 19484 4944 19490 4956
rect 129274 4944 129280 4956
rect 19484 4916 129280 4944
rect 19484 4904 19490 4916
rect 129274 4904 129280 4916
rect 129332 4904 129338 4956
rect 147858 4904 147864 4956
rect 147916 4944 147922 4956
rect 200086 4944 200114 4984
rect 220446 4972 220452 4984
rect 220504 4972 220510 5024
rect 147916 4916 200114 4944
rect 147916 4904 147922 4916
rect 21818 4836 21824 4888
rect 21876 4876 21882 4888
rect 131298 4876 131304 4888
rect 21876 4848 131304 4876
rect 21876 4836 21882 4848
rect 131298 4836 131304 4848
rect 131356 4836 131362 4888
rect 142522 4836 142528 4888
rect 142580 4876 142586 4888
rect 158898 4876 158904 4888
rect 142580 4848 158904 4876
rect 142580 4836 142586 4848
rect 158898 4836 158904 4848
rect 158956 4836 158962 4888
rect 169662 4836 169668 4888
rect 169720 4876 169726 4888
rect 494698 4876 494704 4888
rect 169720 4848 494704 4876
rect 169720 4836 169726 4848
rect 494698 4836 494704 4848
rect 494756 4836 494762 4888
rect 18230 4768 18236 4820
rect 18288 4808 18294 4820
rect 131482 4808 131488 4820
rect 18288 4780 131488 4808
rect 18288 4768 18294 4780
rect 131482 4768 131488 4780
rect 131540 4768 131546 4820
rect 144086 4768 144092 4820
rect 144144 4808 144150 4820
rect 170766 4808 170772 4820
rect 144144 4780 170772 4808
rect 144144 4768 144150 4780
rect 170766 4768 170772 4780
rect 170824 4768 170830 4820
rect 171134 4768 171140 4820
rect 171192 4808 171198 4820
rect 533706 4808 533712 4820
rect 171192 4780 533712 4808
rect 171192 4768 171198 4780
rect 533706 4768 533712 4780
rect 533764 4768 533770 4820
rect 6454 4088 6460 4140
rect 6512 4128 6518 4140
rect 7558 4128 7564 4140
rect 6512 4100 7564 4128
rect 6512 4088 6518 4100
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 140958 4088 140964 4140
rect 141016 4128 141022 4140
rect 144730 4128 144736 4140
rect 141016 4100 144736 4128
rect 141016 4088 141022 4100
rect 144730 4088 144736 4100
rect 144788 4088 144794 4140
rect 148410 4088 148416 4140
rect 148468 4128 148474 4140
rect 153010 4128 153016 4140
rect 148468 4100 153016 4128
rect 148468 4088 148474 4100
rect 153010 4088 153016 4100
rect 153068 4088 153074 4140
rect 225138 4128 225144 4140
rect 156616 4100 225144 4128
rect 125870 4020 125876 4072
rect 125928 4060 125934 4072
rect 139762 4060 139768 4072
rect 125928 4032 139768 4060
rect 125928 4020 125934 4032
rect 139762 4020 139768 4032
rect 139820 4020 139826 4072
rect 147766 4020 147772 4072
rect 147824 4060 147830 4072
rect 156616 4060 156644 4100
rect 225138 4088 225144 4100
rect 225196 4088 225202 4140
rect 343634 4088 343640 4140
rect 343692 4128 343698 4140
rect 351638 4128 351644 4140
rect 343692 4100 351644 4128
rect 343692 4088 343698 4100
rect 351638 4088 351644 4100
rect 351696 4088 351702 4140
rect 352558 4088 352564 4140
rect 352616 4128 352622 4140
rect 355226 4128 355232 4140
rect 352616 4100 355232 4128
rect 352616 4088 352622 4100
rect 355226 4088 355232 4100
rect 355284 4088 355290 4140
rect 357158 4088 357164 4140
rect 357216 4128 357222 4140
rect 367002 4128 367008 4140
rect 357216 4100 367008 4128
rect 357216 4088 357222 4100
rect 367002 4088 367008 4100
rect 367060 4088 367066 4140
rect 389818 4088 389824 4140
rect 389876 4128 389882 4140
rect 394234 4128 394240 4140
rect 389876 4100 394240 4128
rect 389876 4088 389882 4100
rect 394234 4088 394240 4100
rect 394292 4088 394298 4140
rect 147824 4032 156644 4060
rect 147824 4020 147830 4032
rect 156690 4020 156696 4072
rect 156748 4060 156754 4072
rect 228726 4060 228732 4072
rect 156748 4032 228732 4060
rect 156748 4020 156754 4032
rect 228726 4020 228732 4032
rect 228784 4020 228790 4072
rect 303522 4020 303528 4072
rect 303580 4060 303586 4072
rect 310238 4060 310244 4072
rect 303580 4032 310244 4060
rect 303580 4020 303586 4032
rect 310238 4020 310244 4032
rect 310296 4020 310302 4072
rect 344370 4020 344376 4072
rect 344428 4060 344434 4072
rect 358722 4060 358728 4072
rect 344428 4032 358728 4060
rect 344428 4020 344434 4032
rect 358722 4020 358728 4032
rect 358780 4020 358786 4072
rect 373994 4060 374000 4072
rect 364306 4032 374000 4060
rect 86862 3952 86868 4004
rect 86920 3992 86926 4004
rect 137278 3992 137284 4004
rect 86920 3964 137284 3992
rect 86920 3952 86926 3964
rect 137278 3952 137284 3964
rect 137336 3952 137342 4004
rect 149146 3952 149152 4004
rect 149204 3992 149210 4004
rect 239306 3992 239312 4004
rect 149204 3964 239312 3992
rect 149204 3952 149210 3964
rect 239306 3952 239312 3964
rect 239364 3952 239370 4004
rect 251174 3952 251180 4004
rect 251232 3992 251238 4004
rect 252370 3992 252376 4004
rect 251232 3964 252376 3992
rect 251232 3952 251238 3964
rect 252370 3952 252376 3964
rect 252428 3952 252434 4004
rect 307018 3952 307024 4004
rect 307076 3992 307082 4004
rect 318518 3992 318524 4004
rect 307076 3964 318524 3992
rect 307076 3952 307082 3964
rect 318518 3952 318524 3964
rect 318576 3952 318582 4004
rect 322382 3952 322388 4004
rect 322440 3992 322446 4004
rect 329190 3992 329196 4004
rect 322440 3964 329196 3992
rect 322440 3952 322446 3964
rect 329190 3952 329196 3964
rect 329248 3952 329254 4004
rect 353294 3952 353300 4004
rect 353352 3992 353358 4004
rect 364306 3992 364334 4032
rect 373994 4020 374000 4032
rect 374052 4020 374058 4072
rect 370222 3992 370228 4004
rect 353352 3964 364334 3992
rect 367940 3964 370228 3992
rect 353352 3952 353358 3964
rect 69106 3884 69112 3936
rect 69164 3924 69170 3936
rect 135346 3924 135352 3936
rect 69164 3896 135352 3924
rect 69164 3884 69170 3896
rect 135346 3884 135352 3896
rect 135404 3884 135410 3936
rect 150434 3884 150440 3936
rect 150492 3924 150498 3936
rect 258258 3924 258264 3936
rect 150492 3896 258264 3924
rect 150492 3884 150498 3896
rect 258258 3884 258264 3896
rect 258316 3884 258322 3936
rect 276014 3884 276020 3936
rect 276072 3924 276078 3936
rect 276750 3924 276756 3936
rect 276072 3896 276756 3924
rect 276072 3884 276078 3896
rect 276750 3884 276756 3896
rect 276808 3884 276814 3936
rect 317414 3884 317420 3936
rect 317472 3924 317478 3936
rect 330386 3924 330392 3936
rect 317472 3896 330392 3924
rect 317472 3884 317478 3896
rect 330386 3884 330392 3896
rect 330444 3884 330450 3936
rect 333974 3884 333980 3936
rect 334032 3924 334038 3936
rect 340966 3924 340972 3936
rect 334032 3896 340972 3924
rect 334032 3884 334038 3896
rect 340966 3884 340972 3896
rect 341024 3884 341030 3936
rect 342806 3884 342812 3936
rect 342864 3924 342870 3936
rect 367940 3924 367968 3964
rect 370222 3952 370228 3964
rect 370280 3952 370286 4004
rect 370498 3952 370504 4004
rect 370556 3992 370562 4004
rect 378870 3992 378876 4004
rect 370556 3964 378876 3992
rect 370556 3952 370562 3964
rect 378870 3952 378876 3964
rect 378928 3952 378934 4004
rect 342864 3896 367968 3924
rect 342864 3884 342870 3896
rect 369118 3884 369124 3936
rect 369176 3924 369182 3936
rect 372890 3924 372896 3936
rect 369176 3896 372896 3924
rect 369176 3884 369182 3896
rect 372890 3884 372896 3896
rect 372948 3884 372954 3936
rect 62022 3816 62028 3868
rect 62080 3856 62086 3868
rect 128998 3856 129004 3868
rect 62080 3828 129004 3856
rect 62080 3816 62086 3828
rect 128998 3816 129004 3828
rect 129056 3816 129062 3868
rect 144454 3816 144460 3868
rect 144512 3856 144518 3868
rect 160094 3856 160100 3868
rect 144512 3828 160100 3856
rect 144512 3816 144518 3828
rect 160094 3816 160100 3828
rect 160152 3816 160158 3868
rect 166718 3816 166724 3868
rect 166776 3856 166782 3868
rect 458082 3856 458088 3868
rect 166776 3828 458088 3856
rect 166776 3816 166782 3828
rect 458082 3816 458088 3828
rect 458140 3816 458146 3868
rect 461670 3816 461676 3868
rect 461728 3856 461734 3868
rect 471054 3856 471060 3868
rect 461728 3828 471060 3856
rect 461728 3816 461734 3828
rect 471054 3816 471060 3828
rect 471112 3816 471118 3868
rect 9950 3748 9956 3800
rect 10008 3788 10014 3800
rect 88886 3788 88892 3800
rect 10008 3760 88892 3788
rect 10008 3748 10014 3760
rect 88886 3748 88892 3760
rect 88944 3748 88950 3800
rect 93946 3748 93952 3800
rect 94004 3788 94010 3800
rect 137094 3788 137100 3800
rect 94004 3760 137100 3788
rect 94004 3748 94010 3760
rect 137094 3748 137100 3760
rect 137152 3748 137158 3800
rect 143442 3748 143448 3800
rect 143500 3788 143506 3800
rect 151814 3788 151820 3800
rect 143500 3760 151820 3788
rect 143500 3748 143506 3760
rect 151814 3748 151820 3760
rect 151872 3748 151878 3800
rect 176102 3748 176108 3800
rect 176160 3788 176166 3800
rect 472250 3788 472256 3800
rect 176160 3760 472256 3788
rect 176160 3748 176166 3760
rect 472250 3748 472256 3760
rect 472308 3748 472314 3800
rect 39574 3680 39580 3732
rect 39632 3720 39638 3732
rect 129090 3720 129096 3732
rect 39632 3692 129096 3720
rect 39632 3680 39638 3692
rect 129090 3680 129096 3692
rect 129148 3680 129154 3732
rect 140682 3680 140688 3732
rect 140740 3720 140746 3732
rect 161290 3720 161296 3732
rect 140740 3692 161296 3720
rect 140740 3680 140746 3692
rect 161290 3680 161296 3692
rect 161348 3680 161354 3732
rect 177574 3680 177580 3732
rect 177632 3720 177638 3732
rect 480530 3720 480536 3732
rect 177632 3692 480536 3720
rect 177632 3680 177638 3692
rect 480530 3680 480536 3692
rect 480588 3680 480594 3732
rect 17034 3612 17040 3664
rect 17092 3652 17098 3664
rect 131942 3652 131948 3664
rect 17092 3624 131948 3652
rect 17092 3612 17098 3624
rect 131942 3612 131948 3624
rect 132000 3612 132006 3664
rect 143718 3612 143724 3664
rect 143776 3652 143782 3664
rect 167178 3652 167184 3664
rect 143776 3624 167184 3652
rect 143776 3612 143782 3624
rect 167178 3612 167184 3624
rect 167236 3612 167242 3664
rect 177390 3612 177396 3664
rect 177448 3652 177454 3664
rect 181438 3652 181444 3664
rect 177448 3624 181444 3652
rect 177448 3612 177454 3624
rect 181438 3612 181444 3624
rect 181496 3612 181502 3664
rect 185578 3612 185584 3664
rect 185636 3652 185642 3664
rect 487614 3652 487620 3664
rect 185636 3624 487620 3652
rect 185636 3612 185642 3624
rect 487614 3612 487620 3624
rect 487672 3612 487678 3664
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 1728 3556 4384 3584
rect 1728 3544 1734 3556
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 4356 3516 4384 3556
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 10318 3584 10324 3596
rect 5316 3556 10324 3584
rect 5316 3544 5322 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 11974 3584 11980 3596
rect 11112 3556 11980 3584
rect 11112 3544 11118 3556
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 131206 3584 131212 3596
rect 13596 3556 131212 3584
rect 13596 3544 13602 3556
rect 131206 3544 131212 3556
rect 131264 3544 131270 3596
rect 141050 3544 141056 3596
rect 141108 3584 141114 3596
rect 147122 3584 147128 3596
rect 141108 3556 147128 3584
rect 141108 3544 141114 3556
rect 147122 3544 147128 3556
rect 147180 3544 147186 3596
rect 149238 3544 149244 3596
rect 149296 3584 149302 3596
rect 174262 3584 174268 3596
rect 149296 3556 174268 3584
rect 149296 3544 149302 3556
rect 174262 3544 174268 3556
rect 174320 3544 174326 3596
rect 177298 3544 177304 3596
rect 177356 3584 177362 3596
rect 491110 3584 491116 3596
rect 177356 3556 491116 3584
rect 177356 3544 177362 3556
rect 491110 3544 491116 3556
rect 491168 3544 491174 3596
rect 126238 3516 126244 3528
rect 4356 3488 126244 3516
rect 126238 3476 126244 3488
rect 126296 3476 126302 3528
rect 131758 3476 131764 3528
rect 131816 3516 131822 3528
rect 140038 3516 140044 3528
rect 131816 3488 140044 3516
rect 131816 3476 131822 3488
rect 140038 3476 140044 3488
rect 140096 3476 140102 3528
rect 143626 3476 143632 3528
rect 143684 3516 143690 3528
rect 171962 3516 171968 3528
rect 143684 3488 171968 3516
rect 143684 3476 143690 3488
rect 171962 3476 171968 3488
rect 172020 3476 172026 3528
rect 176194 3476 176200 3528
rect 176252 3516 176258 3528
rect 177850 3516 177856 3528
rect 176252 3488 177856 3516
rect 176252 3476 176258 3488
rect 177850 3476 177856 3488
rect 177908 3476 177914 3528
rect 177942 3476 177948 3528
rect 178000 3516 178006 3528
rect 505370 3516 505376 3528
rect 178000 3488 505376 3516
rect 178000 3476 178006 3488
rect 505370 3476 505376 3488
rect 505428 3476 505434 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 507302 3516 507308 3528
rect 506532 3488 507308 3516
rect 506532 3476 506538 3488
rect 507302 3476 507308 3488
rect 507360 3476 507366 3528
rect 531314 3476 531320 3528
rect 531372 3516 531378 3528
rect 532142 3516 532148 3528
rect 531372 3488 532148 3516
rect 531372 3476 531378 3488
rect 532142 3476 532148 3488
rect 532200 3476 532206 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 127618 3448 127624 3460
rect 624 3420 127624 3448
rect 624 3408 630 3420
rect 127618 3408 127624 3420
rect 127676 3408 127682 3460
rect 132954 3408 132960 3460
rect 133012 3448 133018 3460
rect 140130 3448 140136 3460
rect 133012 3420 140136 3448
rect 133012 3408 133018 3420
rect 140130 3408 140136 3420
rect 140188 3408 140194 3460
rect 144546 3408 144552 3460
rect 144604 3448 144610 3460
rect 175458 3448 175464 3460
rect 144604 3420 175464 3448
rect 144604 3408 144610 3420
rect 175458 3408 175464 3420
rect 175516 3408 175522 3460
rect 177758 3408 177764 3460
rect 177816 3448 177822 3460
rect 508866 3448 508872 3460
rect 177816 3420 508872 3448
rect 177816 3408 177822 3420
rect 508866 3408 508872 3420
rect 508924 3408 508930 3460
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 147674 3340 147680 3392
rect 147732 3380 147738 3392
rect 156690 3380 156696 3392
rect 147732 3352 156696 3380
rect 147732 3340 147738 3352
rect 156690 3340 156696 3352
rect 156748 3340 156754 3392
rect 189718 3380 189724 3392
rect 161446 3352 189724 3380
rect 141510 3272 141516 3324
rect 141568 3312 141574 3324
rect 143534 3312 143540 3324
rect 141568 3284 143540 3312
rect 141568 3272 141574 3284
rect 143534 3272 143540 3284
rect 143592 3272 143598 3324
rect 147214 3204 147220 3256
rect 147272 3244 147278 3256
rect 161446 3244 161474 3352
rect 189718 3340 189724 3352
rect 189776 3340 189782 3392
rect 218054 3340 218060 3392
rect 218112 3380 218118 3392
rect 219250 3380 219256 3392
rect 218112 3352 219256 3380
rect 218112 3340 218118 3352
rect 219250 3340 219256 3352
rect 219308 3340 219314 3392
rect 242894 3340 242900 3392
rect 242952 3380 242958 3392
rect 244090 3380 244096 3392
rect 242952 3352 244096 3380
rect 242952 3340 242958 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 302142 3340 302148 3392
rect 302200 3380 302206 3392
rect 309042 3380 309048 3392
rect 302200 3352 309048 3380
rect 302200 3340 302206 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 322290 3340 322296 3392
rect 322348 3380 322354 3392
rect 325602 3380 325608 3392
rect 322348 3352 325608 3380
rect 322348 3340 322354 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 329098 3340 329104 3392
rect 329156 3380 329162 3392
rect 336274 3380 336280 3392
rect 329156 3352 336280 3380
rect 329156 3340 329162 3352
rect 336274 3340 336280 3352
rect 336332 3340 336338 3392
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 374086 3340 374092 3392
rect 374144 3380 374150 3392
rect 375282 3380 375288 3392
rect 374144 3352 375288 3380
rect 374144 3340 374150 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382366 3340 382372 3392
rect 382424 3380 382430 3392
rect 383562 3380 383568 3392
rect 382424 3352 383568 3380
rect 382424 3340 382430 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 390646 3340 390652 3392
rect 390704 3380 390710 3392
rect 391842 3380 391848 3392
rect 390704 3352 391848 3380
rect 390704 3340 390710 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 431954 3340 431960 3392
rect 432012 3380 432018 3392
rect 433242 3380 433248 3392
rect 432012 3352 433248 3380
rect 432012 3340 432018 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 465718 3340 465724 3392
rect 465776 3380 465782 3392
rect 469858 3380 469864 3392
rect 465776 3352 469864 3380
rect 465776 3340 465782 3352
rect 469858 3340 469864 3352
rect 469916 3340 469922 3392
rect 175918 3272 175924 3324
rect 175976 3312 175982 3324
rect 177942 3312 177948 3324
rect 175976 3284 177948 3312
rect 175976 3272 175982 3284
rect 177942 3272 177948 3284
rect 178000 3272 178006 3324
rect 186130 3312 186136 3324
rect 178052 3284 186136 3312
rect 147272 3216 161474 3244
rect 147272 3204 147278 3216
rect 171870 3204 171876 3256
rect 171928 3244 171934 3256
rect 176654 3244 176660 3256
rect 171928 3216 176660 3244
rect 171928 3204 171934 3216
rect 176654 3204 176660 3216
rect 176712 3204 176718 3256
rect 142246 3136 142252 3188
rect 142304 3176 142310 3188
rect 150618 3176 150624 3188
rect 142304 3148 150624 3176
rect 142304 3136 142310 3148
rect 150618 3136 150624 3148
rect 150676 3136 150682 3188
rect 172054 3068 172060 3120
rect 172112 3108 172118 3120
rect 178052 3108 178080 3284
rect 186130 3272 186136 3284
rect 186188 3272 186194 3324
rect 319806 3272 319812 3324
rect 319864 3312 319870 3324
rect 322106 3312 322112 3324
rect 319864 3284 322112 3312
rect 319864 3272 319870 3284
rect 322106 3272 322112 3284
rect 322164 3272 322170 3324
rect 334066 3272 334072 3324
rect 334124 3312 334130 3324
rect 337470 3312 337476 3324
rect 334124 3284 337476 3312
rect 334124 3272 334130 3284
rect 337470 3272 337476 3284
rect 337528 3272 337534 3324
rect 322198 3204 322204 3256
rect 322256 3244 322262 3256
rect 326798 3244 326804 3256
rect 322256 3216 326804 3244
rect 322256 3204 322262 3216
rect 326798 3204 326804 3216
rect 326856 3204 326862 3256
rect 384390 3204 384396 3256
rect 384448 3244 384454 3256
rect 387150 3244 387156 3256
rect 384448 3216 387156 3244
rect 384448 3204 384454 3216
rect 387150 3204 387156 3216
rect 387208 3204 387214 3256
rect 309226 3136 309232 3188
rect 309284 3176 309290 3188
rect 317322 3176 317328 3188
rect 309284 3148 317328 3176
rect 309284 3136 309290 3148
rect 317322 3136 317328 3148
rect 317380 3136 317386 3188
rect 482278 3136 482284 3188
rect 482336 3176 482342 3188
rect 485222 3176 485228 3188
rect 482336 3148 485228 3176
rect 482336 3136 482342 3148
rect 485222 3136 485228 3148
rect 485280 3136 485286 3188
rect 172112 3080 178080 3108
rect 172112 3068 172118 3080
rect 327074 3068 327080 3120
rect 327132 3108 327138 3120
rect 331582 3108 331588 3120
rect 327132 3080 331588 3108
rect 327132 3068 327138 3080
rect 331582 3068 331588 3080
rect 331640 3068 331646 3120
rect 347038 3068 347044 3120
rect 347096 3108 347102 3120
rect 354030 3108 354036 3120
rect 347096 3080 354036 3108
rect 347096 3068 347102 3080
rect 354030 3068 354036 3080
rect 354088 3068 354094 3120
rect 140038 3000 140044 3052
rect 140096 3040 140102 3052
rect 141142 3040 141148 3052
rect 140096 3012 141148 3040
rect 140096 3000 140102 3012
rect 141142 3000 141148 3012
rect 141200 3000 141206 3052
rect 145558 3000 145564 3052
rect 145616 3040 145622 3052
rect 154206 3040 154212 3052
rect 145616 3012 154212 3040
rect 145616 3000 145622 3012
rect 154206 3000 154212 3012
rect 154264 3000 154270 3052
rect 175550 3000 175556 3052
rect 175608 3040 175614 3052
rect 185578 3040 185584 3052
rect 175608 3012 185584 3040
rect 175608 3000 175614 3012
rect 185578 3000 185584 3012
rect 185636 3000 185642 3052
rect 330478 3000 330484 3052
rect 330536 3040 330542 3052
rect 333882 3040 333888 3052
rect 330536 3012 333888 3040
rect 330536 3000 330542 3012
rect 333882 3000 333888 3012
rect 333940 3000 333946 3052
rect 362954 3000 362960 3052
rect 363012 3040 363018 3052
rect 365806 3040 365812 3052
rect 363012 3012 365812 3040
rect 363012 3000 363018 3012
rect 365806 3000 365812 3012
rect 365864 3000 365870 3052
rect 308398 2932 308404 2984
rect 308456 2972 308462 2984
rect 311434 2972 311440 2984
rect 308456 2944 311440 2972
rect 308456 2932 308462 2944
rect 311434 2932 311440 2944
rect 311492 2932 311498 2984
rect 407114 1776 407120 1828
rect 407172 1816 407178 1828
rect 408402 1816 408408 1828
rect 407172 1788 408408 1816
rect 407172 1776 407178 1788
rect 408402 1776 408408 1788
rect 408460 1776 408466 1828
rect 415394 1776 415400 1828
rect 415452 1816 415458 1828
rect 416682 1816 416688 1828
rect 415452 1788 416688 1816
rect 415452 1776 415458 1788
rect 416682 1776 416688 1788
rect 416740 1776 416746 1828
rect 440234 1776 440240 1828
rect 440292 1816 440298 1828
rect 441522 1816 441528 1828
rect 440292 1788 441528 1816
rect 440292 1776 440298 1788
rect 441522 1776 441528 1788
rect 441580 1776 441586 1828
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 207664 700680 207716 700732
rect 218980 700680 219032 700732
rect 192484 700612 192536 700664
rect 267648 700612 267700 700664
rect 206284 700544 206336 700596
rect 283840 700544 283892 700596
rect 203524 700476 203576 700528
rect 348792 700476 348844 700528
rect 200764 700408 200816 700460
rect 413652 700408 413704 700460
rect 199384 700340 199436 700392
rect 478512 700340 478564 700392
rect 137836 700272 137888 700324
rect 190460 700272 190512 700324
rect 198004 700272 198056 700324
rect 543464 700272 543516 700324
rect 105452 699660 105504 699712
rect 106924 699660 106976 699712
rect 193864 699660 193916 699712
rect 202788 699660 202840 699712
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 196624 683136 196676 683188
rect 580172 683136 580224 683188
rect 3424 656888 3476 656940
rect 116584 656888 116636 656940
rect 3424 632068 3476 632120
rect 7564 632068 7616 632120
rect 193956 630640 194008 630692
rect 580172 630640 580224 630692
rect 120724 616836 120776 616888
rect 580172 616836 580224 616888
rect 3332 579640 3384 579692
rect 17224 579640 17276 579692
rect 194048 576852 194100 576904
rect 579620 576852 579672 576904
rect 120816 563048 120868 563100
rect 580172 563048 580224 563100
rect 3332 553392 3384 553444
rect 116676 553392 116728 553444
rect 3332 527824 3384 527876
rect 8944 527824 8996 527876
rect 194140 524424 194192 524476
rect 579804 524424 579856 524476
rect 3332 514768 3384 514820
rect 190552 514768 190604 514820
rect 120908 510620 120960 510672
rect 579988 510620 580040 510672
rect 118700 485052 118752 485104
rect 580540 485052 580592 485104
rect 221464 470568 221516 470620
rect 579620 470568 579672 470620
rect 3056 462340 3108 462392
rect 189724 462340 189776 462392
rect 3884 461592 3936 461644
rect 48964 461592 49016 461644
rect 121000 456764 121052 456816
rect 579620 456764 579672 456816
rect 2964 448536 3016 448588
rect 84844 448536 84896 448588
rect 3332 422288 3384 422340
rect 10324 422288 10376 422340
rect 192576 418140 192628 418192
rect 579712 418140 579764 418192
rect 3332 409844 3384 409896
rect 189080 409844 189132 409896
rect 118608 404336 118660 404388
rect 580172 404336 580224 404388
rect 3332 397468 3384 397520
rect 112444 397468 112496 397520
rect 3332 371220 3384 371272
rect 84936 371220 84988 371272
rect 360844 364352 360896 364404
rect 580172 364352 580224 364404
rect 118516 351908 118568 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 121092 345040 121144 345092
rect 3148 318792 3200 318844
rect 13084 318792 13136 318844
rect 359464 311856 359516 311908
rect 580172 311856 580224 311908
rect 3332 304988 3384 305040
rect 185584 304988 185636 305040
rect 146944 298120 146996 298172
rect 580172 298120 580224 298172
rect 3240 266364 3292 266416
rect 18604 266364 18656 266416
rect 202144 258068 202196 258120
rect 580172 258068 580224 258120
rect 2872 253920 2924 253972
rect 190644 253920 190696 253972
rect 122104 244264 122156 244316
rect 580172 244264 580224 244316
rect 194232 231820 194284 231872
rect 579804 231820 579856 231872
rect 225604 218016 225656 218068
rect 579988 218016 580040 218068
rect 3332 213936 3384 213988
rect 31024 213936 31076 213988
rect 147036 205640 147088 205692
rect 580172 205640 580224 205692
rect 3332 201492 3384 201544
rect 189264 201492 189316 201544
rect 192668 191836 192720 191888
rect 580172 191836 580224 191888
rect 3332 187688 3384 187740
rect 119344 187688 119396 187740
rect 224224 178032 224276 178084
rect 580172 178032 580224 178084
rect 122196 165588 122248 165640
rect 580172 165588 580224 165640
rect 3332 162868 3384 162920
rect 14464 162868 14516 162920
rect 3792 160692 3844 160744
rect 189356 160692 189408 160744
rect 192760 151784 192812 151836
rect 579988 151784 580040 151836
rect 3516 149880 3568 149932
rect 3792 149880 3844 149932
rect 3516 148316 3568 148368
rect 191196 148316 191248 148368
rect 119252 146956 119304 147008
rect 234620 146956 234672 147008
rect 3608 146888 3660 146940
rect 190828 146888 190880 146940
rect 118976 145596 119028 145648
rect 299480 145596 299532 145648
rect 3792 145528 3844 145580
rect 189448 145528 189500 145580
rect 23480 144236 23532 144288
rect 189540 144236 189592 144288
rect 119068 144168 119120 144220
rect 364340 144168 364392 144220
rect 118240 142944 118292 142996
rect 146944 142944 146996 142996
rect 3884 142876 3936 142928
rect 191104 142876 191156 142928
rect 119160 142808 119212 142860
rect 429200 142808 429252 142860
rect 118424 141516 118476 141568
rect 147036 141516 147088 141568
rect 88340 141448 88392 141500
rect 191012 141448 191064 141500
rect 118884 141380 118936 141432
rect 494060 141380 494112 141432
rect 185584 140496 185636 140548
rect 192024 140496 192076 140548
rect 153200 140156 153252 140208
rect 190920 140156 190972 140208
rect 118056 140088 118108 140140
rect 169760 140088 169812 140140
rect 118792 140020 118844 140072
rect 558920 140020 558972 140072
rect 118148 139544 118200 139596
rect 122104 139544 122156 139596
rect 118332 139476 118384 139528
rect 122196 139476 122248 139528
rect 3608 139408 3660 139460
rect 191932 139408 191984 139460
rect 7656 136688 7708 136740
rect 117320 136688 117372 136740
rect 3516 136620 3568 136672
rect 119436 136620 119488 136672
rect 9036 135260 9088 135312
rect 117320 135260 117372 135312
rect 21364 133900 21416 133952
rect 117320 133900 117372 133952
rect 14464 133832 14516 133884
rect 117412 133832 117464 133884
rect 31024 132404 31076 132456
rect 117320 132404 117372 132456
rect 18604 131044 18656 131096
rect 117320 131044 117372 131096
rect 189172 129752 189224 129804
rect 189632 129752 189684 129804
rect 13084 129684 13136 129736
rect 117320 129684 117372 129736
rect 84936 128256 84988 128308
rect 117320 128256 117372 128308
rect 10324 126896 10376 126948
rect 117320 126896 117372 126948
rect 189264 126896 189316 126948
rect 189632 126896 189684 126948
rect 48964 124108 49016 124160
rect 117320 124108 117372 124160
rect 8944 122748 8996 122800
rect 117320 122748 117372 122800
rect 17224 121388 17276 121440
rect 117320 121388 117372 121440
rect 189080 121388 189132 121440
rect 189356 121388 189408 121440
rect 7564 120028 7616 120080
rect 117320 120028 117372 120080
rect 4804 118600 4856 118652
rect 117320 118600 117372 118652
rect 40040 117240 40092 117292
rect 117320 117240 117372 117292
rect 106924 115880 106976 115932
rect 117320 115880 117372 115932
rect 189724 111800 189776 111852
rect 580080 111800 580132 111852
rect 3332 111732 3384 111784
rect 21364 111732 21416 111784
rect 191932 108944 191984 108996
rect 207664 108944 207716 108996
rect 191932 107584 191984 107636
rect 206284 107584 206336 107636
rect 191932 106224 191984 106276
rect 203524 106224 203576 106276
rect 193128 104796 193180 104848
rect 200764 104796 200816 104848
rect 193128 102484 193180 102536
rect 199384 102484 199436 102536
rect 191932 101124 191984 101176
rect 198004 101124 198056 101176
rect 192392 100648 192444 100700
rect 196624 100648 196676 100700
rect 192116 98472 192168 98524
rect 193956 98472 194008 98524
rect 192208 97452 192260 97504
rect 194048 97452 194100 97504
rect 191932 96432 191984 96484
rect 194140 96432 194192 96484
rect 193128 95140 193180 95192
rect 221464 95140 221516 95192
rect 360936 94528 360988 94580
rect 580172 94528 580224 94580
rect 359556 94460 359608 94512
rect 579988 94460 580040 94512
rect 193128 92420 193180 92472
rect 360844 92420 360896 92472
rect 193128 90992 193180 91044
rect 359464 90992 359516 91044
rect 193128 89632 193180 89684
rect 202144 89632 202196 89684
rect 192944 88952 192996 89004
rect 225604 88952 225656 89004
rect 193036 87592 193088 87644
rect 224224 87592 224276 87644
rect 580172 86368 580224 86420
rect 580816 86368 580868 86420
rect 193128 85484 193180 85536
rect 360936 85484 360988 85536
rect 3332 84192 3384 84244
rect 120632 84192 120684 84244
rect 193128 84124 193180 84176
rect 359556 84124 359608 84176
rect 189080 80724 189132 80776
rect 580264 80724 580316 80776
rect 188988 80656 189040 80708
rect 580356 80656 580408 80708
rect 193128 80112 193180 80164
rect 526444 80112 526496 80164
rect 3700 79976 3752 80028
rect 127072 79976 127124 80028
rect 127256 79976 127308 80028
rect 130200 79976 130252 80028
rect 127164 79908 127216 79960
rect 129924 79908 129976 79960
rect 130798 79908 130850 79960
rect 130982 79908 131034 79960
rect 131534 79908 131586 79960
rect 121092 79840 121144 79892
rect 129464 79840 129516 79892
rect 129556 79840 129608 79892
rect 131258 79840 131310 79892
rect 126888 79772 126940 79824
rect 131166 79772 131218 79824
rect 131028 79704 131080 79756
rect 131350 79772 131402 79824
rect 126336 79636 126388 79688
rect 119436 79568 119488 79620
rect 127624 79568 127676 79620
rect 131120 79636 131172 79688
rect 131994 79908 132046 79960
rect 131718 79840 131770 79892
rect 131902 79840 131954 79892
rect 131856 79704 131908 79756
rect 132270 79840 132322 79892
rect 132822 79840 132874 79892
rect 131948 79636 132000 79688
rect 132224 79568 132276 79620
rect 132546 79772 132598 79824
rect 133374 79908 133426 79960
rect 133558 79908 133610 79960
rect 133742 79908 133794 79960
rect 133834 79908 133886 79960
rect 133190 79840 133242 79892
rect 133696 79772 133748 79824
rect 133512 79704 133564 79756
rect 132592 79636 132644 79688
rect 132684 79636 132736 79688
rect 132868 79636 132920 79688
rect 133328 79636 133380 79688
rect 133788 79636 133840 79688
rect 132500 79568 132552 79620
rect 134202 79908 134254 79960
rect 135214 79908 135266 79960
rect 134662 79840 134714 79892
rect 134938 79840 134990 79892
rect 135122 79840 135174 79892
rect 134064 79636 134116 79688
rect 134800 79636 134852 79688
rect 135076 79636 135128 79688
rect 135168 79636 135220 79688
rect 135628 79636 135680 79688
rect 135858 79840 135910 79892
rect 135950 79840 136002 79892
rect 134156 79568 134208 79620
rect 120632 79500 120684 79552
rect 129372 79500 129424 79552
rect 129464 79500 129516 79552
rect 135904 79568 135956 79620
rect 135444 79500 135496 79552
rect 136686 79908 136738 79960
rect 136778 79908 136830 79960
rect 136870 79908 136922 79960
rect 137514 79908 137566 79960
rect 138158 79908 138210 79960
rect 136594 79840 136646 79892
rect 136824 79772 136876 79824
rect 136732 79704 136784 79756
rect 136548 79636 136600 79688
rect 116676 79432 116728 79484
rect 127624 79432 127676 79484
rect 135352 79432 135404 79484
rect 136272 79432 136324 79484
rect 137882 79840 137934 79892
rect 137100 79636 137152 79688
rect 138020 79636 138072 79688
rect 138894 79840 138946 79892
rect 139078 79840 139130 79892
rect 139538 79908 139590 79960
rect 139262 79840 139314 79892
rect 138296 79636 138348 79688
rect 138480 79636 138532 79688
rect 139124 79636 139176 79688
rect 139722 79840 139774 79892
rect 139584 79636 139636 79688
rect 139216 79568 139268 79620
rect 139814 79772 139866 79824
rect 137008 79500 137060 79552
rect 139400 79500 139452 79552
rect 137744 79432 137796 79484
rect 139768 79432 139820 79484
rect 140366 79908 140418 79960
rect 140458 79908 140510 79960
rect 140550 79908 140602 79960
rect 140090 79840 140142 79892
rect 140182 79840 140234 79892
rect 140320 79772 140372 79824
rect 140412 79704 140464 79756
rect 140642 79840 140694 79892
rect 141010 79840 141062 79892
rect 140228 79636 140280 79688
rect 140044 79568 140096 79620
rect 141378 79908 141430 79960
rect 141470 79908 141522 79960
rect 141240 79636 141292 79688
rect 140780 79568 140832 79620
rect 141148 79568 141200 79620
rect 140504 79500 140556 79552
rect 141056 79500 141108 79552
rect 141746 79908 141798 79960
rect 141838 79908 141890 79960
rect 141930 79908 141982 79960
rect 142022 79908 142074 79960
rect 142114 79908 142166 79960
rect 142298 79908 142350 79960
rect 142758 79908 142810 79960
rect 142942 79908 142994 79960
rect 143034 79908 143086 79960
rect 141700 79772 141752 79824
rect 141884 79636 141936 79688
rect 140780 79432 140832 79484
rect 141792 79432 141844 79484
rect 142390 79840 142442 79892
rect 142482 79840 142534 79892
rect 142574 79840 142626 79892
rect 142344 79704 142396 79756
rect 142068 79636 142120 79688
rect 142252 79636 142304 79688
rect 143586 79840 143638 79892
rect 142988 79772 143040 79824
rect 143770 79908 143822 79960
rect 143724 79772 143776 79824
rect 143632 79704 143684 79756
rect 142712 79636 142764 79688
rect 142896 79636 142948 79688
rect 143448 79636 143500 79688
rect 143540 79636 143592 79688
rect 143954 79840 144006 79892
rect 142436 79500 142488 79552
rect 144782 79908 144834 79960
rect 144874 79908 144926 79960
rect 144414 79840 144466 79892
rect 144506 79840 144558 79892
rect 143908 79568 143960 79620
rect 144736 79772 144788 79824
rect 144828 79772 144880 79824
rect 144644 79568 144696 79620
rect 144092 79500 144144 79552
rect 142896 79432 142948 79484
rect 144368 79432 144420 79484
rect 145242 79908 145294 79960
rect 145518 79908 145570 79960
rect 145058 79772 145110 79824
rect 145288 79500 145340 79552
rect 145196 79432 145248 79484
rect 146162 79840 146214 79892
rect 146254 79840 146306 79892
rect 146346 79840 146398 79892
rect 146208 79636 146260 79688
rect 145656 79500 145708 79552
rect 146990 79908 147042 79960
rect 147174 79908 147226 79960
rect 146622 79840 146674 79892
rect 146806 79840 146858 79892
rect 146760 79500 146812 79552
rect 145932 79432 145984 79484
rect 146300 79432 146352 79484
rect 146944 79636 146996 79688
rect 144920 79364 144972 79416
rect 145104 79364 145156 79416
rect 145840 79364 145892 79416
rect 146484 79364 146536 79416
rect 147266 79840 147318 79892
rect 147358 79840 147410 79892
rect 147542 79772 147594 79824
rect 147404 79704 147456 79756
rect 147220 79636 147272 79688
rect 147496 79636 147548 79688
rect 147128 79568 147180 79620
rect 147910 79908 147962 79960
rect 148186 79908 148238 79960
rect 148278 79908 148330 79960
rect 148370 79908 148422 79960
rect 148738 79908 148790 79960
rect 149382 79908 149434 79960
rect 149934 79908 149986 79960
rect 150026 79908 150078 79960
rect 147818 79840 147870 79892
rect 147726 79772 147778 79824
rect 147772 79636 147824 79688
rect 148554 79840 148606 79892
rect 148324 79704 148376 79756
rect 148232 79636 148284 79688
rect 148416 79636 148468 79688
rect 148922 79840 148974 79892
rect 149014 79840 149066 79892
rect 149198 79840 149250 79892
rect 148784 79772 148836 79824
rect 148876 79704 148928 79756
rect 149152 79704 149204 79756
rect 149428 79636 149480 79688
rect 149658 79840 149710 79892
rect 148600 79568 148652 79620
rect 148692 79568 148744 79620
rect 150210 79840 150262 79892
rect 150394 79840 150446 79892
rect 150486 79840 150538 79892
rect 150670 79840 150722 79892
rect 149980 79704 150032 79756
rect 149888 79636 149940 79688
rect 150256 79636 150308 79688
rect 150578 79772 150630 79824
rect 150716 79704 150768 79756
rect 150624 79636 150676 79688
rect 150164 79500 150216 79552
rect 149244 79432 149296 79484
rect 149520 79432 149572 79484
rect 148968 79364 149020 79416
rect 149336 79364 149388 79416
rect 149796 79364 149848 79416
rect 150440 79500 150492 79552
rect 151130 79908 151182 79960
rect 151314 79908 151366 79960
rect 151406 79908 151458 79960
rect 151498 79908 151550 79960
rect 151958 79908 152010 79960
rect 152510 79908 152562 79960
rect 152602 79908 152654 79960
rect 152786 79908 152838 79960
rect 152970 79908 153022 79960
rect 153062 79908 153114 79960
rect 153154 79908 153206 79960
rect 153246 79908 153298 79960
rect 151038 79840 151090 79892
rect 151222 79840 151274 79892
rect 151084 79704 151136 79756
rect 151176 79704 151228 79756
rect 151268 79704 151320 79756
rect 151360 79636 151412 79688
rect 151774 79840 151826 79892
rect 151866 79840 151918 79892
rect 151728 79636 151780 79688
rect 151912 79636 151964 79688
rect 150900 79568 150952 79620
rect 151452 79568 151504 79620
rect 151636 79568 151688 79620
rect 151820 79568 151872 79620
rect 152234 79840 152286 79892
rect 152418 79840 152470 79892
rect 152142 79772 152194 79824
rect 152280 79704 152332 79756
rect 152372 79704 152424 79756
rect 152648 79704 152700 79756
rect 152832 79704 152884 79756
rect 153108 79704 153160 79756
rect 152556 79568 152608 79620
rect 152188 79500 152240 79552
rect 153292 79636 153344 79688
rect 153200 79500 153252 79552
rect 153016 79432 153068 79484
rect 153522 79772 153574 79824
rect 153614 79772 153666 79824
rect 153568 79636 153620 79688
rect 153890 79908 153942 79960
rect 153982 79908 154034 79960
rect 154074 79908 154126 79960
rect 154166 79908 154218 79960
rect 154258 79908 154310 79960
rect 154350 79908 154402 79960
rect 154028 79704 154080 79756
rect 153844 79636 153896 79688
rect 153936 79568 153988 79620
rect 154534 79908 154586 79960
rect 154626 79908 154678 79960
rect 154718 79908 154770 79960
rect 154994 79908 155046 79960
rect 155086 79908 155138 79960
rect 155178 79908 155230 79960
rect 155270 79908 155322 79960
rect 154304 79704 154356 79756
rect 154396 79704 154448 79756
rect 154672 79704 154724 79756
rect 154488 79636 154540 79688
rect 154580 79568 154632 79620
rect 155132 79772 155184 79824
rect 154948 79704 155000 79756
rect 155040 79568 155092 79620
rect 153752 79500 153804 79552
rect 155224 79500 155276 79552
rect 155454 79908 155506 79960
rect 155408 79704 155460 79756
rect 156098 79908 156150 79960
rect 156190 79908 156242 79960
rect 156282 79908 156334 79960
rect 155730 79840 155782 79892
rect 155914 79840 155966 79892
rect 156006 79840 156058 79892
rect 155684 79636 155736 79688
rect 155868 79704 155920 79756
rect 156374 79840 156426 79892
rect 156236 79704 156288 79756
rect 156144 79568 156196 79620
rect 156328 79568 156380 79620
rect 156558 79840 156610 79892
rect 156834 79908 156886 79960
rect 157110 79908 157162 79960
rect 157202 79908 157254 79960
rect 157386 79908 157438 79960
rect 157478 79908 157530 79960
rect 157570 79908 157622 79960
rect 157662 79908 157714 79960
rect 156788 79772 156840 79824
rect 156512 79568 156564 79620
rect 155776 79500 155828 79552
rect 156420 79500 156472 79552
rect 156604 79500 156656 79552
rect 157294 79840 157346 79892
rect 157156 79704 157208 79756
rect 157248 79636 157300 79688
rect 157340 79568 157392 79620
rect 157846 79840 157898 79892
rect 157616 79636 157668 79688
rect 157524 79568 157576 79620
rect 157064 79500 157116 79552
rect 157800 79568 157852 79620
rect 158306 79908 158358 79960
rect 158398 79908 158450 79960
rect 158582 79908 158634 79960
rect 158674 79908 158726 79960
rect 159134 79908 159186 79960
rect 159226 79908 159278 79960
rect 159502 79908 159554 79960
rect 159686 79908 159738 79960
rect 159778 79908 159830 79960
rect 160054 79908 160106 79960
rect 160146 79908 160198 79960
rect 160238 79908 160290 79960
rect 160422 79908 160474 79960
rect 160606 79908 160658 79960
rect 160790 79908 160842 79960
rect 160882 79908 160934 79960
rect 161250 79908 161302 79960
rect 161434 79908 161486 79960
rect 161710 79908 161762 79960
rect 162078 79908 162130 79960
rect 158030 79840 158082 79892
rect 158214 79840 158266 79892
rect 158122 79772 158174 79824
rect 158352 79772 158404 79824
rect 158444 79772 158496 79824
rect 158582 79772 158634 79824
rect 158260 79704 158312 79756
rect 158858 79840 158910 79892
rect 158950 79840 159002 79892
rect 158168 79636 158220 79688
rect 158628 79636 158680 79688
rect 157984 79500 158036 79552
rect 159180 79636 159232 79688
rect 158996 79568 159048 79620
rect 159088 79568 159140 79620
rect 158904 79500 158956 79552
rect 159272 79500 159324 79552
rect 159548 79568 159600 79620
rect 159824 79568 159876 79620
rect 154212 79432 154264 79484
rect 158352 79432 158404 79484
rect 158628 79432 158680 79484
rect 160330 79840 160382 79892
rect 160192 79636 160244 79688
rect 160468 79772 160520 79824
rect 160560 79704 160612 79756
rect 160744 79636 160796 79688
rect 160836 79568 160888 79620
rect 161066 79840 161118 79892
rect 161158 79840 161210 79892
rect 161296 79704 161348 79756
rect 160284 79500 160336 79552
rect 160468 79500 160520 79552
rect 160928 79500 160980 79552
rect 161112 79500 161164 79552
rect 161894 79840 161946 79892
rect 161802 79772 161854 79824
rect 161664 79704 161716 79756
rect 162262 79772 162314 79824
rect 162216 79568 162268 79620
rect 161572 79500 161624 79552
rect 162032 79500 162084 79552
rect 161480 79432 161532 79484
rect 162538 79908 162590 79960
rect 162814 79908 162866 79960
rect 162906 79908 162958 79960
rect 162400 79636 162452 79688
rect 162814 79772 162866 79824
rect 162492 79432 162544 79484
rect 162768 79432 162820 79484
rect 162998 79772 163050 79824
rect 163826 79908 163878 79960
rect 163918 79908 163970 79960
rect 163458 79840 163510 79892
rect 163550 79840 163602 79892
rect 163734 79840 163786 79892
rect 163504 79704 163556 79756
rect 163596 79636 163648 79688
rect 163688 79636 163740 79688
rect 164010 79772 164062 79824
rect 164470 79908 164522 79960
rect 164286 79840 164338 79892
rect 164562 79840 164614 79892
rect 163964 79636 164016 79688
rect 164332 79704 164384 79756
rect 163780 79568 163832 79620
rect 163872 79568 163924 79620
rect 164056 79568 164108 79620
rect 164240 79568 164292 79620
rect 165758 79908 165810 79960
rect 164930 79840 164982 79892
rect 165022 79840 165074 79892
rect 165114 79840 165166 79892
rect 165298 79840 165350 79892
rect 165666 79840 165718 79892
rect 164976 79704 165028 79756
rect 165574 79772 165626 79824
rect 165160 79704 165212 79756
rect 165252 79704 165304 79756
rect 165712 79704 165764 79756
rect 165942 79908 165994 79960
rect 166034 79908 166086 79960
rect 166126 79908 166178 79960
rect 165068 79636 165120 79688
rect 165528 79636 165580 79688
rect 165804 79636 165856 79688
rect 166402 79840 166454 79892
rect 165988 79772 166040 79824
rect 166080 79772 166132 79824
rect 166218 79772 166270 79824
rect 166172 79636 166224 79688
rect 165988 79568 166040 79620
rect 164424 79500 164476 79552
rect 164700 79500 164752 79552
rect 163044 79432 163096 79484
rect 163504 79432 163556 79484
rect 152648 79364 152700 79416
rect 3976 79296 4028 79348
rect 130200 79228 130252 79280
rect 132684 79228 132736 79280
rect 134524 79228 134576 79280
rect 140136 79228 140188 79280
rect 129372 79160 129424 79212
rect 140044 79160 140096 79212
rect 137284 79092 137336 79144
rect 140136 79092 140188 79144
rect 140964 79296 141016 79348
rect 141976 79296 142028 79348
rect 149244 79296 149296 79348
rect 158076 79364 158128 79416
rect 158536 79364 158588 79416
rect 165620 79364 165672 79416
rect 165896 79364 165948 79416
rect 166356 79432 166408 79484
rect 166862 79908 166914 79960
rect 166770 79840 166822 79892
rect 166954 79840 167006 79892
rect 166816 79568 166868 79620
rect 166632 79500 166684 79552
rect 167138 79908 167190 79960
rect 167598 79908 167650 79960
rect 167230 79840 167282 79892
rect 167414 79840 167466 79892
rect 167782 79908 167834 79960
rect 167874 79908 167926 79960
rect 167966 79908 168018 79960
rect 168058 79908 168110 79960
rect 167092 79704 167144 79756
rect 167184 79704 167236 79756
rect 167460 79704 167512 79756
rect 167552 79636 167604 79688
rect 167920 79704 167972 79756
rect 167736 79568 167788 79620
rect 167828 79568 167880 79620
rect 168794 79908 168846 79960
rect 169438 79908 169490 79960
rect 168610 79840 168662 79892
rect 168656 79704 168708 79756
rect 168288 79568 168340 79620
rect 166908 79432 166960 79484
rect 168104 79432 168156 79484
rect 168886 79840 168938 79892
rect 169346 79840 169398 79892
rect 169530 79840 169582 79892
rect 169024 79568 169076 79620
rect 168840 79500 168892 79552
rect 169392 79704 169444 79756
rect 169484 79636 169536 79688
rect 169806 79908 169858 79960
rect 169898 79908 169950 79960
rect 169990 79908 170042 79960
rect 170174 79908 170226 79960
rect 170818 79908 170870 79960
rect 171554 79908 171606 79960
rect 171646 79908 171698 79960
rect 169760 79704 169812 79756
rect 169300 79568 169352 79620
rect 170450 79840 170502 79892
rect 170542 79840 170594 79892
rect 170128 79704 170180 79756
rect 170496 79704 170548 79756
rect 170036 79636 170088 79688
rect 170036 79500 170088 79552
rect 170680 79636 170732 79688
rect 171370 79840 171422 79892
rect 171324 79704 171376 79756
rect 171600 79636 171652 79688
rect 171232 79500 171284 79552
rect 171830 79908 171882 79960
rect 171922 79908 171974 79960
rect 172014 79908 172066 79960
rect 172474 79908 172526 79960
rect 172566 79908 172618 79960
rect 172750 79908 172802 79960
rect 172934 79908 172986 79960
rect 173118 79908 173170 79960
rect 171784 79704 171836 79756
rect 166632 79364 166684 79416
rect 167000 79364 167052 79416
rect 167276 79364 167328 79416
rect 168564 79364 168616 79416
rect 169576 79296 169628 79348
rect 170312 79432 170364 79484
rect 171416 79432 171468 79484
rect 172198 79840 172250 79892
rect 172014 79772 172066 79824
rect 172106 79772 172158 79824
rect 172060 79568 172112 79620
rect 172290 79772 172342 79824
rect 172152 79500 172204 79552
rect 172244 79432 172296 79484
rect 170128 79364 170180 79416
rect 170496 79364 170548 79416
rect 172336 79364 172388 79416
rect 172612 79500 172664 79552
rect 173302 79840 173354 79892
rect 173026 79772 173078 79824
rect 172704 79432 172756 79484
rect 172980 79636 173032 79688
rect 173486 79908 173538 79960
rect 173578 79908 173630 79960
rect 173670 79908 173722 79960
rect 173854 79908 173906 79960
rect 173578 79772 173630 79824
rect 173532 79636 173584 79688
rect 173624 79636 173676 79688
rect 173440 79568 173492 79620
rect 173256 79500 173308 79552
rect 173716 79500 173768 79552
rect 174222 79908 174274 79960
rect 174314 79908 174366 79960
rect 174406 79908 174458 79960
rect 174498 79908 174550 79960
rect 174590 79908 174642 79960
rect 174774 79908 174826 79960
rect 174866 79908 174918 79960
rect 175050 79908 175102 79960
rect 175326 79908 175378 79960
rect 175970 79908 176022 79960
rect 176154 79908 176206 79960
rect 176338 79908 176390 79960
rect 176522 79908 176574 79960
rect 176614 79908 176666 79960
rect 176706 79908 176758 79960
rect 176798 79908 176850 79960
rect 176890 79908 176942 79960
rect 176982 79908 177034 79960
rect 177074 79908 177126 79960
rect 174084 79500 174136 79552
rect 174452 79704 174504 79756
rect 174774 79772 174826 79824
rect 175142 79840 175194 79892
rect 175096 79704 175148 79756
rect 175188 79704 175240 79756
rect 176062 79840 176114 79892
rect 176016 79704 176068 79756
rect 176108 79704 176160 79756
rect 174544 79568 174596 79620
rect 174452 79500 174504 79552
rect 174544 79432 174596 79484
rect 174728 79500 174780 79552
rect 175372 79636 175424 79688
rect 172796 79364 172848 79416
rect 173164 79364 173216 79416
rect 175464 79364 175516 79416
rect 176476 79704 176528 79756
rect 176568 79704 176620 79756
rect 176384 79636 176436 79688
rect 176844 79704 176896 79756
rect 176936 79704 176988 79756
rect 176844 79500 176896 79552
rect 177258 79908 177310 79960
rect 177350 79908 177402 79960
rect 188896 80044 188948 80096
rect 580448 80044 580500 80096
rect 177442 79840 177494 79892
rect 177718 79840 177770 79892
rect 177304 79772 177356 79824
rect 177212 79704 177264 79756
rect 177810 79772 177862 79824
rect 178454 79908 178506 79960
rect 178914 79908 178966 79960
rect 179972 79976 180024 80028
rect 179696 79908 179748 79960
rect 179282 79840 179334 79892
rect 179788 79840 179840 79892
rect 180248 79772 180300 79824
rect 194232 79772 194284 79824
rect 180524 79704 180576 79756
rect 181720 79568 181772 79620
rect 177396 79432 177448 79484
rect 178040 79432 178092 79484
rect 178132 79432 178184 79484
rect 415400 79500 415452 79552
rect 189724 79364 189776 79416
rect 173072 79296 173124 79348
rect 176752 79296 176804 79348
rect 177120 79296 177172 79348
rect 179972 79296 180024 79348
rect 140964 79160 141016 79212
rect 141884 79160 141936 79212
rect 144460 79160 144512 79212
rect 173348 79228 173400 79280
rect 175004 79228 175056 79280
rect 176384 79228 176436 79280
rect 179880 79228 179932 79280
rect 157432 79160 157484 79212
rect 159364 79160 159416 79212
rect 160100 79160 160152 79212
rect 158076 79092 158128 79144
rect 164056 79092 164108 79144
rect 112444 79024 112496 79076
rect 130016 78956 130068 79008
rect 130844 78956 130896 79008
rect 84844 78888 84896 78940
rect 140044 78888 140096 78940
rect 144460 78888 144512 78940
rect 144920 78888 144972 78940
rect 129372 78820 129424 78872
rect 134156 78820 134208 78872
rect 135352 78820 135404 78872
rect 155316 78888 155368 78940
rect 158352 78956 158404 79008
rect 160100 78956 160152 79008
rect 162584 78956 162636 79008
rect 162860 78956 162912 79008
rect 163228 78956 163280 79008
rect 163596 78956 163648 79008
rect 164516 79024 164568 79076
rect 164884 79024 164936 79076
rect 165804 79160 165856 79212
rect 176292 79160 176344 79212
rect 177304 79160 177356 79212
rect 527180 79296 527232 79348
rect 180524 79228 180576 79280
rect 192484 79228 192536 79280
rect 181720 79160 181772 79212
rect 193864 79160 193916 79212
rect 166540 79092 166592 79144
rect 171784 79092 171836 79144
rect 172428 79092 172480 79144
rect 175280 79092 175332 79144
rect 168564 79024 168616 79076
rect 169576 79024 169628 79076
rect 178868 79092 178920 79144
rect 176660 79024 176712 79076
rect 178132 79024 178184 79076
rect 179880 79024 179932 79076
rect 192668 79092 192720 79144
rect 170128 78888 170180 78940
rect 122104 78616 122156 78668
rect 133880 78752 133932 78804
rect 135996 78752 136048 78804
rect 136180 78752 136232 78804
rect 154212 78820 154264 78872
rect 130844 78684 130896 78736
rect 138572 78684 138624 78736
rect 139216 78684 139268 78736
rect 140044 78684 140096 78736
rect 140504 78684 140556 78736
rect 144368 78616 144420 78668
rect 155224 78684 155276 78736
rect 158812 78820 158864 78872
rect 172888 78888 172940 78940
rect 173164 78888 173216 78940
rect 176200 78956 176252 79008
rect 192760 78956 192812 79008
rect 178592 78888 178644 78940
rect 177856 78820 177908 78872
rect 178040 78820 178092 78872
rect 180524 78820 180576 78872
rect 158536 78752 158588 78804
rect 162400 78752 162452 78804
rect 164792 78752 164844 78804
rect 169576 78752 169628 78804
rect 170128 78752 170180 78804
rect 178408 78752 178460 78804
rect 157340 78684 157392 78736
rect 161112 78684 161164 78736
rect 161204 78684 161256 78736
rect 162584 78684 162636 78736
rect 162676 78684 162728 78736
rect 167184 78684 167236 78736
rect 167460 78684 167512 78736
rect 161020 78616 161072 78668
rect 162400 78616 162452 78668
rect 164240 78616 164292 78668
rect 164424 78616 164476 78668
rect 164608 78616 164660 78668
rect 164792 78616 164844 78668
rect 166172 78616 166224 78668
rect 170128 78616 170180 78668
rect 150716 78548 150768 78600
rect 177764 78684 177816 78736
rect 171600 78616 171652 78668
rect 174820 78616 174872 78668
rect 175832 78616 175884 78668
rect 177212 78616 177264 78668
rect 177396 78616 177448 78668
rect 173072 78548 173124 78600
rect 178776 78548 178828 78600
rect 580632 78548 580684 78600
rect 134432 78480 134484 78532
rect 134800 78480 134852 78532
rect 136364 78480 136416 78532
rect 137192 78480 137244 78532
rect 146576 78480 146628 78532
rect 171048 78480 171100 78532
rect 172888 78480 172940 78532
rect 173808 78480 173860 78532
rect 175648 78480 175700 78532
rect 176568 78480 176620 78532
rect 176752 78480 176804 78532
rect 179144 78480 179196 78532
rect 180248 78480 180300 78532
rect 188896 78480 188948 78532
rect 130660 78412 130712 78464
rect 138664 78412 138716 78464
rect 140136 78412 140188 78464
rect 154580 78412 154632 78464
rect 161572 78412 161624 78464
rect 162032 78412 162084 78464
rect 164056 78412 164108 78464
rect 171508 78412 171560 78464
rect 158720 78344 158772 78396
rect 163964 78344 164016 78396
rect 170128 78344 170180 78396
rect 454040 78412 454092 78464
rect 171784 78344 171836 78396
rect 460940 78344 460992 78396
rect 129464 78276 129516 78328
rect 139584 78276 139636 78328
rect 140136 78276 140188 78328
rect 140872 78276 140924 78328
rect 161388 78276 161440 78328
rect 166172 78276 166224 78328
rect 167368 78276 167420 78328
rect 467840 78276 467892 78328
rect 127716 78208 127768 78260
rect 134524 78208 134576 78260
rect 161664 78208 161716 78260
rect 162676 78208 162728 78260
rect 167552 78208 167604 78260
rect 474740 78208 474792 78260
rect 118700 78140 118752 78192
rect 139400 78140 139452 78192
rect 157800 78140 157852 78192
rect 164608 78140 164660 78192
rect 172612 78140 172664 78192
rect 172980 78140 173032 78192
rect 175372 78140 175424 78192
rect 96620 78072 96672 78124
rect 138020 78072 138072 78124
rect 145472 78072 145524 78124
rect 147312 78072 147364 78124
rect 150808 78072 150860 78124
rect 78680 78004 78732 78056
rect 136824 78004 136876 78056
rect 145196 78004 145248 78056
rect 159916 78072 159968 78124
rect 165804 78072 165856 78124
rect 170312 78072 170364 78124
rect 10324 77936 10376 77988
rect 129556 77936 129608 77988
rect 131488 77936 131540 77988
rect 132408 77936 132460 77988
rect 145380 77936 145432 77988
rect 147588 77936 147640 77988
rect 131672 77868 131724 77920
rect 131948 77868 132000 77920
rect 129004 77800 129056 77852
rect 135260 77800 135312 77852
rect 129188 77732 129240 77784
rect 139032 77732 139084 77784
rect 128360 77664 128412 77716
rect 140780 77664 140832 77716
rect 172704 78004 172756 78056
rect 172980 78004 173032 78056
rect 173992 78004 174044 78056
rect 174452 78004 174504 78056
rect 175740 78072 175792 78124
rect 179880 78140 179932 78192
rect 557540 78140 557592 78192
rect 175832 78004 175884 78056
rect 574100 78072 574152 78124
rect 581000 78004 581052 78056
rect 162860 77936 162912 77988
rect 162216 77868 162268 77920
rect 173440 77936 173492 77988
rect 175924 77936 175976 77988
rect 176476 77936 176528 77988
rect 187884 77936 187936 77988
rect 168196 77732 168248 77784
rect 176200 77868 176252 77920
rect 177212 77868 177264 77920
rect 582380 77936 582432 77988
rect 171508 77800 171560 77852
rect 177304 77800 177356 77852
rect 187884 77800 187936 77852
rect 580172 77868 580224 77920
rect 176384 77732 176436 77784
rect 129832 77596 129884 77648
rect 136732 77596 136784 77648
rect 148048 77596 148100 77648
rect 148416 77596 148468 77648
rect 169576 77664 169628 77716
rect 177212 77664 177264 77716
rect 172428 77596 172480 77648
rect 174820 77596 174872 77648
rect 178776 77596 178828 77648
rect 130752 77528 130804 77580
rect 132132 77528 132184 77580
rect 135260 77528 135312 77580
rect 140872 77528 140924 77580
rect 147956 77528 148008 77580
rect 148232 77528 148284 77580
rect 148692 77528 148744 77580
rect 172336 77528 172388 77580
rect 180616 77528 180668 77580
rect 190460 77528 190512 77580
rect 131856 77460 131908 77512
rect 135628 77460 135680 77512
rect 156144 77460 156196 77512
rect 168288 77460 168340 77512
rect 171048 77460 171100 77512
rect 177488 77460 177540 77512
rect 129280 77392 129332 77444
rect 132040 77392 132092 77444
rect 132132 77392 132184 77444
rect 133144 77392 133196 77444
rect 140688 77392 140740 77444
rect 143172 77392 143224 77444
rect 143724 77392 143776 77444
rect 144368 77392 144420 77444
rect 157892 77392 157944 77444
rect 158812 77392 158864 77444
rect 160376 77392 160428 77444
rect 165436 77392 165488 77444
rect 168380 77392 168432 77444
rect 173808 77392 173860 77444
rect 130384 77324 130436 77376
rect 137836 77324 137888 77376
rect 164332 77324 164384 77376
rect 177672 77324 177724 77376
rect 126244 77256 126296 77308
rect 130568 77256 130620 77308
rect 132408 77256 132460 77308
rect 134248 77256 134300 77308
rect 134524 77256 134576 77308
rect 136456 77256 136508 77308
rect 163688 77256 163740 77308
rect 165344 77256 165396 77308
rect 165804 77256 165856 77308
rect 166632 77256 166684 77308
rect 178224 77256 178276 77308
rect 179788 77256 179840 77308
rect 126980 77188 127032 77240
rect 140412 77188 140464 77240
rect 144828 77188 144880 77240
rect 185032 77188 185084 77240
rect 104900 76984 104952 77036
rect 145104 77120 145156 77172
rect 145748 77120 145800 77172
rect 146208 77120 146260 77172
rect 147680 77120 147732 77172
rect 147772 77120 147824 77172
rect 148048 77120 148100 77172
rect 173072 77120 173124 77172
rect 173624 77120 173676 77172
rect 175280 77120 175332 77172
rect 233240 77120 233292 77172
rect 155408 77052 155460 77104
rect 222936 77052 222988 77104
rect 138848 76984 138900 77036
rect 150624 76984 150676 77036
rect 150900 76984 150952 77036
rect 168196 76984 168248 77036
rect 259460 76984 259512 77036
rect 91100 76916 91152 76968
rect 137652 76916 137704 76968
rect 145380 76916 145432 76968
rect 146116 76916 146168 76968
rect 153292 76916 153344 76968
rect 153752 76916 153804 76968
rect 159364 76916 159416 76968
rect 273536 76916 273588 76968
rect 85580 76848 85632 76900
rect 136364 76848 136416 76900
rect 151452 76848 151504 76900
rect 267740 76848 267792 76900
rect 84200 76780 84252 76832
rect 136640 76780 136692 76832
rect 160284 76780 160336 76832
rect 280344 76780 280396 76832
rect 67640 76712 67692 76764
rect 131856 76712 131908 76764
rect 142344 76712 142396 76764
rect 143080 76712 143132 76764
rect 160652 76712 160704 76764
rect 311900 76712 311952 76764
rect 59360 76644 59412 76696
rect 135168 76644 135220 76696
rect 158904 76644 158956 76696
rect 336740 76644 336792 76696
rect 34520 76576 34572 76628
rect 11060 76508 11112 76560
rect 127164 76508 127216 76560
rect 133052 76576 133104 76628
rect 133512 76576 133564 76628
rect 142160 76576 142212 76628
rect 142620 76576 142672 76628
rect 142712 76576 142764 76628
rect 142896 76576 142948 76628
rect 147680 76576 147732 76628
rect 148508 76576 148560 76628
rect 160284 76576 160336 76628
rect 160744 76576 160796 76628
rect 172796 76576 172848 76628
rect 173164 76576 173216 76628
rect 177856 76576 177908 76628
rect 361580 76576 361632 76628
rect 132684 76508 132736 76560
rect 133696 76508 133748 76560
rect 147128 76508 147180 76560
rect 148140 76508 148192 76560
rect 149612 76508 149664 76560
rect 150072 76508 150124 76560
rect 161848 76508 161900 76560
rect 398840 76508 398892 76560
rect 133236 76440 133288 76492
rect 156696 76440 156748 76492
rect 178500 76440 178552 76492
rect 131488 76372 131540 76424
rect 132224 76372 132276 76424
rect 145472 76372 145524 76424
rect 146024 76372 146076 76424
rect 149612 76372 149664 76424
rect 149888 76372 149940 76424
rect 156420 76372 156472 76424
rect 143816 76304 143868 76356
rect 144092 76304 144144 76356
rect 164608 76304 164660 76356
rect 165252 76304 165304 76356
rect 146392 76236 146444 76288
rect 149888 76236 149940 76288
rect 153384 76236 153436 76288
rect 153568 76236 153620 76288
rect 169852 76236 169904 76288
rect 170312 76236 170364 76288
rect 172704 76372 172756 76424
rect 173348 76372 173400 76424
rect 172796 76304 172848 76356
rect 173532 76304 173584 76356
rect 179144 76236 179196 76288
rect 153292 76168 153344 76220
rect 153844 76168 153896 76220
rect 168472 76168 168524 76220
rect 175648 76168 175700 76220
rect 146392 76100 146444 76152
rect 147220 76100 147272 76152
rect 157524 76100 157576 76152
rect 179052 76100 179104 76152
rect 160376 76032 160428 76084
rect 160560 76032 160612 76084
rect 168656 76032 168708 76084
rect 170956 76032 171008 76084
rect 171508 76032 171560 76084
rect 172152 76032 172204 76084
rect 141424 75964 141476 76016
rect 141608 75964 141660 76016
rect 150624 75964 150676 76016
rect 151360 75964 151412 76016
rect 152004 75964 152056 76016
rect 152740 75964 152792 76016
rect 153016 75964 153068 76016
rect 153936 75964 153988 76016
rect 167000 75964 167052 76016
rect 176016 75964 176068 76016
rect 129096 75896 129148 75948
rect 133604 75896 133656 75948
rect 138020 75896 138072 75948
rect 141332 75896 141384 75948
rect 149060 75896 149112 75948
rect 149244 75896 149296 75948
rect 150808 75896 150860 75948
rect 151176 75896 151228 75948
rect 151728 75896 151780 75948
rect 152464 75896 152516 75948
rect 153200 75896 153252 75948
rect 154212 75896 154264 75948
rect 155040 75896 155092 75948
rect 158536 75896 158588 75948
rect 159732 75896 159784 75948
rect 159916 75896 159968 75948
rect 166540 75896 166592 75948
rect 166724 75896 166776 75948
rect 168472 75896 168524 75948
rect 168932 75896 168984 75948
rect 169116 75896 169168 75948
rect 169668 75896 169720 75948
rect 170312 75896 170364 75948
rect 170772 75896 170824 75948
rect 171140 75896 171192 75948
rect 171692 75896 171744 75948
rect 118516 75828 118568 75880
rect 580908 75828 580960 75880
rect 141332 75760 141384 75812
rect 141792 75760 141844 75812
rect 145932 75760 145984 75812
rect 191840 75760 191892 75812
rect 280344 75760 280396 75812
rect 283196 75760 283248 75812
rect 148968 75692 149020 75744
rect 220820 75692 220872 75744
rect 144644 75624 144696 75676
rect 176200 75624 176252 75676
rect 177764 75624 177816 75676
rect 256700 75624 256752 75676
rect 131304 75556 131356 75608
rect 136180 75556 136232 75608
rect 153200 75556 153252 75608
rect 154028 75556 154080 75608
rect 157708 75556 157760 75608
rect 159732 75556 159784 75608
rect 159824 75556 159876 75608
rect 262864 75556 262916 75608
rect 130936 75488 130988 75540
rect 140596 75488 140648 75540
rect 151912 75488 151964 75540
rect 274640 75488 274692 75540
rect 311900 75488 311952 75540
rect 320548 75488 320600 75540
rect 127072 75420 127124 75472
rect 140320 75420 140372 75472
rect 169208 75420 169260 75472
rect 114560 75352 114612 75404
rect 139124 75352 139176 75404
rect 159180 75352 159232 75404
rect 137284 75284 137336 75336
rect 157708 75284 157760 75336
rect 164332 75284 164384 75336
rect 165068 75284 165120 75336
rect 75920 75216 75972 75268
rect 131304 75216 131356 75268
rect 134248 75216 134300 75268
rect 134708 75216 134760 75268
rect 135628 75216 135680 75268
rect 136272 75216 136324 75268
rect 138388 75216 138440 75268
rect 139308 75216 139360 75268
rect 139584 75216 139636 75268
rect 140228 75216 140280 75268
rect 155316 75216 155368 75268
rect 156880 75216 156932 75268
rect 161664 75216 161716 75268
rect 161848 75216 161900 75268
rect 163136 75216 163188 75268
rect 163504 75216 163556 75268
rect 164516 75216 164568 75268
rect 164884 75216 164936 75268
rect 53840 75148 53892 75200
rect 134340 75148 134392 75200
rect 135076 75148 135128 75200
rect 135720 75148 135772 75200
rect 136548 75148 136600 75200
rect 162860 75148 162912 75200
rect 163228 75148 163280 75200
rect 164608 75148 164660 75200
rect 164976 75148 165028 75200
rect 131304 75080 131356 75132
rect 132500 75080 132552 75132
rect 163136 75080 163188 75132
rect 163780 75080 163832 75132
rect 164240 75080 164292 75132
rect 165160 75080 165212 75132
rect 166172 75352 166224 75404
rect 166540 75352 166592 75404
rect 171140 75352 171192 75404
rect 172060 75352 172112 75404
rect 173808 75420 173860 75472
rect 485780 75420 485832 75472
rect 496820 75352 496872 75404
rect 165896 75284 165948 75336
rect 166448 75284 166500 75336
rect 169392 75284 169444 75336
rect 499580 75284 499632 75336
rect 165620 75216 165672 75268
rect 166172 75216 166224 75268
rect 167000 75216 167052 75268
rect 167828 75216 167880 75268
rect 170588 75216 170640 75268
rect 514760 75216 514812 75268
rect 165804 75148 165856 75200
rect 166264 75148 166316 75200
rect 175096 75148 175148 75200
rect 175924 75148 175976 75200
rect 543740 75148 543792 75200
rect 173900 75080 173952 75132
rect 174452 75080 174504 75132
rect 134892 75012 134944 75064
rect 160192 75012 160244 75064
rect 160652 75012 160704 75064
rect 161572 75012 161624 75064
rect 162124 75012 162176 75064
rect 163228 75012 163280 75064
rect 163872 75012 163924 75064
rect 178132 75012 178184 75064
rect 179236 75012 179288 75064
rect 142528 74944 142580 74996
rect 142988 74944 143040 74996
rect 165160 74944 165212 74996
rect 165436 74944 165488 74996
rect 160284 74740 160336 74792
rect 160928 74740 160980 74792
rect 143816 74672 143868 74724
rect 144184 74672 144236 74724
rect 168564 74672 168616 74724
rect 169484 74672 169536 74724
rect 148600 74468 148652 74520
rect 230480 74468 230532 74520
rect 157616 74400 157668 74452
rect 242808 74400 242860 74452
rect 155500 74332 155552 74384
rect 248972 74332 249024 74384
rect 93860 74264 93912 74316
rect 137928 74264 137980 74316
rect 150164 74264 150216 74316
rect 244372 74264 244424 74316
rect 89720 74196 89772 74248
rect 137560 74196 137612 74248
rect 157616 74196 157668 74248
rect 256792 74196 256844 74248
rect 86960 74128 87012 74180
rect 137468 74128 137520 74180
rect 154672 74128 154724 74180
rect 261484 74128 261536 74180
rect 57980 74060 58032 74112
rect 134984 74060 135036 74112
rect 161112 74060 161164 74112
rect 282184 74060 282236 74112
rect 51080 73992 51132 74044
rect 134616 73992 134668 74044
rect 151912 73992 151964 74044
rect 152556 73992 152608 74044
rect 157064 73992 157116 74044
rect 281816 73992 281868 74044
rect 41420 73924 41472 73976
rect 133788 73924 133840 73976
rect 158444 73924 158496 73976
rect 290464 73924 290516 73976
rect 31760 73856 31812 73908
rect 132132 73856 132184 73908
rect 155868 73856 155920 73908
rect 295984 73856 296036 73908
rect 177304 73788 177356 73840
rect 177672 73788 177724 73840
rect 178776 73788 178828 73840
rect 446404 73788 446456 73840
rect 157616 73720 157668 73772
rect 226524 73720 226576 73772
rect 132776 73652 132828 73704
rect 133420 73652 133472 73704
rect 156236 73652 156288 73704
rect 226432 73652 226484 73704
rect 158168 73584 158220 73636
rect 178040 73584 178092 73636
rect 169024 73516 169076 73568
rect 177304 73516 177356 73568
rect 170496 73448 170548 73500
rect 177764 73448 177816 73500
rect 127624 73176 127676 73228
rect 130292 73176 130344 73228
rect 136824 73176 136876 73228
rect 141516 73176 141568 73228
rect 176108 73108 176160 73160
rect 580172 73108 580224 73160
rect 156328 73040 156380 73092
rect 255320 73040 255372 73092
rect 71780 72632 71832 72684
rect 135996 72972 136048 73024
rect 175096 72972 175148 73024
rect 281356 72972 281408 73024
rect 130936 72904 130988 72956
rect 159732 72904 159784 72956
rect 281448 72904 281500 72956
rect 130200 72700 130252 72752
rect 159548 72836 159600 72888
rect 282000 72836 282052 72888
rect 159456 72768 159508 72820
rect 281908 72768 281960 72820
rect 295340 72768 295392 72820
rect 300308 72768 300360 72820
rect 158996 72700 159048 72752
rect 299388 72700 299440 72752
rect 129832 72632 129884 72684
rect 130476 72632 130528 72684
rect 158352 72632 158404 72684
rect 311164 72632 311216 72684
rect 102140 72564 102192 72616
rect 138940 72564 138992 72616
rect 165252 72564 165304 72616
rect 347780 72564 347832 72616
rect 82820 72496 82872 72548
rect 137744 72496 137796 72548
rect 159272 72496 159324 72548
rect 349068 72496 349120 72548
rect 143172 72428 143224 72480
rect 155960 72428 156012 72480
rect 167276 72428 167328 72480
rect 417424 72428 417476 72480
rect 168380 72360 168432 72412
rect 264980 72360 265032 72412
rect 178500 72292 178552 72344
rect 275284 72292 275336 72344
rect 159088 72224 159140 72276
rect 244280 72224 244332 72276
rect 135444 71748 135496 71800
rect 141884 71748 141936 71800
rect 273536 71748 273588 71800
rect 276020 71748 276072 71800
rect 283196 71680 283248 71732
rect 289360 71680 289412 71732
rect 3424 71612 3476 71664
rect 9036 71612 9088 71664
rect 179144 71612 179196 71664
rect 195244 71612 195296 71664
rect 255320 71612 255372 71664
rect 297364 71612 297416 71664
rect 154764 71544 154816 71596
rect 257344 71544 257396 71596
rect 155224 71476 155276 71528
rect 260196 71476 260248 71528
rect 155040 71408 155092 71460
rect 272524 71408 272576 71460
rect 272892 71408 272944 71460
rect 284300 71408 284352 71460
rect 156604 71340 156656 71392
rect 280988 71340 281040 71392
rect 158904 71272 158956 71324
rect 305736 71272 305788 71324
rect 318156 71272 318208 71324
rect 332600 71272 332652 71324
rect 144736 71204 144788 71256
rect 178316 71204 178368 71256
rect 179052 71204 179104 71256
rect 334716 71204 334768 71256
rect 159916 71136 159968 71188
rect 345664 71136 345716 71188
rect 167552 71068 167604 71120
rect 456064 71068 456116 71120
rect 110420 71000 110472 71052
rect 138572 71000 138624 71052
rect 167736 71000 167788 71052
rect 467104 71000 467156 71052
rect 178040 70320 178092 70372
rect 230848 70320 230900 70372
rect 156052 70252 156104 70304
rect 226340 70252 226392 70304
rect 130844 70184 130896 70236
rect 202328 70184 202380 70236
rect 226432 70184 226484 70236
rect 273996 70184 274048 70236
rect 158536 70116 158588 70168
rect 254584 70116 254636 70168
rect 256792 70116 256844 70168
rect 280804 70116 280856 70168
rect 156972 70048 157024 70100
rect 263048 70048 263100 70100
rect 310244 70048 310296 70100
rect 312544 70048 312596 70100
rect 157708 69980 157760 70032
rect 265624 69980 265676 70032
rect 155776 69912 155828 69964
rect 271144 69912 271196 69964
rect 281356 69912 281408 69964
rect 285772 69912 285824 69964
rect 299388 69912 299440 69964
rect 309784 69912 309836 69964
rect 3424 69844 3476 69896
rect 190736 69844 190788 69896
rect 244280 69844 244332 69896
rect 349804 69844 349856 69896
rect 165344 69776 165396 69828
rect 425060 69776 425112 69828
rect 446404 69776 446456 69828
rect 460296 69776 460348 69828
rect 170404 69708 170456 69760
rect 512000 69708 512052 69760
rect 2780 69640 2832 69692
rect 130016 69640 130068 69692
rect 176476 69640 176528 69692
rect 539600 69640 539652 69692
rect 178040 69572 178092 69624
rect 178316 69572 178368 69624
rect 178868 69572 178920 69624
rect 224960 69572 225012 69624
rect 226524 69572 226576 69624
rect 274088 69572 274140 69624
rect 179420 69504 179472 69556
rect 211068 69504 211120 69556
rect 310428 69504 310480 69556
rect 318248 69504 318300 69556
rect 154672 69436 154724 69488
rect 181996 69436 182048 69488
rect 281908 69232 281960 69284
rect 284392 69232 284444 69284
rect 445484 69232 445536 69284
rect 447140 69232 447192 69284
rect 282000 69164 282052 69216
rect 284484 69164 284536 69216
rect 195244 68960 195296 69012
rect 201132 68960 201184 69012
rect 281448 68960 281500 69012
rect 298744 68960 298796 69012
rect 336740 68960 336792 69012
rect 339500 68960 339552 69012
rect 222936 68892 222988 68944
rect 294604 68892 294656 68944
rect 145564 68824 145616 68876
rect 193220 68824 193272 68876
rect 242808 68824 242860 68876
rect 318064 68824 318116 68876
rect 156880 68756 156932 68808
rect 269856 68756 269908 68808
rect 281816 68756 281868 68808
rect 316684 68756 316736 68808
rect 178960 68688 179012 68740
rect 300400 68688 300452 68740
rect 332600 68688 332652 68740
rect 340144 68688 340196 68740
rect 159640 68620 159692 68672
rect 303160 68620 303212 68672
rect 320548 68620 320600 68672
rect 359556 68620 359608 68672
rect 167092 68552 167144 68604
rect 407120 68552 407172 68604
rect 167184 68484 167236 68536
rect 420184 68484 420236 68536
rect 167276 68416 167328 68468
rect 460204 68416 460256 68468
rect 169208 68348 169260 68400
rect 498200 68348 498252 68400
rect 170312 68280 170364 68332
rect 514852 68280 514904 68332
rect 289360 68212 289412 68264
rect 300492 68212 300544 68264
rect 142804 67532 142856 67584
rect 145564 67532 145616 67584
rect 262864 67532 262916 67584
rect 267004 67532 267056 67584
rect 248972 67328 249024 67380
rect 259552 67328 259604 67380
rect 264980 67328 265032 67380
rect 273444 67328 273496 67380
rect 226340 67260 226392 67312
rect 279424 67260 279476 67312
rect 211068 67192 211120 67244
rect 269120 67192 269172 67244
rect 230848 67124 230900 67176
rect 318156 67124 318208 67176
rect 181996 67056 182048 67108
rect 285680 67056 285732 67108
rect 158260 66988 158312 67040
rect 271604 66988 271656 67040
rect 276020 66988 276072 67040
rect 282276 66988 282328 67040
rect 284300 66988 284352 67040
rect 302976 66988 303028 67040
rect 224960 66920 225012 66972
rect 348700 66920 348752 66972
rect 2872 66852 2924 66904
rect 129924 66852 129976 66904
rect 164792 66852 164844 66904
rect 437480 66852 437532 66904
rect 201132 66172 201184 66224
rect 203524 66172 203576 66224
rect 260196 66172 260248 66224
rect 263508 66172 263560 66224
rect 407120 66172 407172 66224
rect 410524 66172 410576 66224
rect 447140 66172 447192 66224
rect 450636 66172 450688 66224
rect 202328 66104 202380 66156
rect 205364 66104 205416 66156
rect 339500 65764 339552 65816
rect 345756 65764 345808 65816
rect 284392 65628 284444 65680
rect 300124 65628 300176 65680
rect 284484 65560 284536 65612
rect 300216 65560 300268 65612
rect 349068 65560 349120 65612
rect 359464 65560 359516 65612
rect 164700 65492 164752 65544
rect 434720 65492 434772 65544
rect 285772 64880 285824 64932
rect 289084 64880 289136 64932
rect 294604 64336 294656 64388
rect 301504 64336 301556 64388
rect 417424 64336 417476 64388
rect 422944 64336 422996 64388
rect 285680 64268 285732 64320
rect 294052 64268 294104 64320
rect 160652 64200 160704 64252
rect 380900 64200 380952 64252
rect 174636 64132 174688 64184
rect 568580 64132 568632 64184
rect 282276 64064 282328 64116
rect 289360 64064 289412 64116
rect 254584 63996 254636 64048
rect 260472 63996 260524 64048
rect 269120 63860 269172 63912
rect 271880 63860 271932 63912
rect 263048 63724 263100 63776
rect 265440 63724 265492 63776
rect 259552 63520 259604 63572
rect 263416 63520 263468 63572
rect 282184 63452 282236 63504
rect 287888 63452 287940 63504
rect 300400 63112 300452 63164
rect 307668 63112 307720 63164
rect 300492 63044 300544 63096
rect 303712 63044 303764 63096
rect 280988 62908 281040 62960
rect 302332 62908 302384 62960
rect 261484 62840 261536 62892
rect 276664 62840 276716 62892
rect 280896 62840 280948 62892
rect 302240 62840 302292 62892
rect 460296 62840 460348 62892
rect 464344 62840 464396 62892
rect 145472 62772 145524 62824
rect 197360 62772 197412 62824
rect 261576 62772 261628 62824
rect 284300 62772 284352 62824
rect 348700 62772 348752 62824
rect 351920 62772 351972 62824
rect 439504 62772 439556 62824
rect 463792 62772 463844 62824
rect 124220 62092 124272 62144
rect 127716 62092 127768 62144
rect 297364 62092 297416 62144
rect 302884 62092 302936 62144
rect 475384 62092 475436 62144
rect 479524 62092 479576 62144
rect 271604 62024 271656 62076
rect 277952 62024 278004 62076
rect 280804 62024 280856 62076
rect 287704 62024 287756 62076
rect 311164 61888 311216 61940
rect 315304 61888 315356 61940
rect 340144 61684 340196 61736
rect 344284 61684 344336 61736
rect 359556 61412 359608 61464
rect 361672 61412 361724 61464
rect 7564 61344 7616 61396
rect 130108 61344 130160 61396
rect 301504 61344 301556 61396
rect 313924 61344 313976 61396
rect 318248 61344 318300 61396
rect 334624 61344 334676 61396
rect 289360 60800 289412 60852
rect 291936 60800 291988 60852
rect 192576 60664 192628 60716
rect 580172 60664 580224 60716
rect 265440 60596 265492 60648
rect 269764 60596 269816 60648
rect 269856 60596 269908 60648
rect 274732 60596 274784 60648
rect 142712 60460 142764 60512
rect 148416 60460 148468 60512
rect 289176 60324 289228 60376
rect 293960 60324 294012 60376
rect 312544 60256 312596 60308
rect 315396 60256 315448 60308
rect 148324 60188 148376 60240
rect 223580 60188 223632 60240
rect 257344 60188 257396 60240
rect 261484 60188 261536 60240
rect 294052 60188 294104 60240
rect 303068 60188 303120 60240
rect 303712 60188 303764 60240
rect 326344 60188 326396 60240
rect 450636 60188 450688 60240
rect 458824 60188 458876 60240
rect 168840 60120 168892 60172
rect 491300 60120 491352 60172
rect 171876 60052 171928 60104
rect 529940 60052 529992 60104
rect 117320 59984 117372 60036
rect 129464 59984 129516 60036
rect 174544 59984 174596 60036
rect 564440 59984 564492 60036
rect 302240 59712 302292 59764
rect 306012 59712 306064 59764
rect 287888 59644 287940 59696
rect 290556 59644 290608 59696
rect 302332 59576 302384 59628
rect 306104 59576 306156 59628
rect 463792 59372 463844 59424
rect 467196 59372 467248 59424
rect 205364 59304 205416 59356
rect 210424 59304 210476 59356
rect 260472 59304 260524 59356
rect 262220 59304 262272 59356
rect 263508 59304 263560 59356
rect 268844 59304 268896 59356
rect 303252 59304 303304 59356
rect 305828 59304 305880 59356
rect 334716 59304 334768 59356
rect 337384 59304 337436 59356
rect 272524 58896 272576 58948
rect 280988 58896 281040 58948
rect 271880 58828 271932 58880
rect 286416 58828 286468 58880
rect 144184 58760 144236 58812
rect 171876 58760 171928 58812
rect 273444 58760 273496 58812
rect 283748 58760 283800 58812
rect 284300 58760 284352 58812
rect 301320 58760 301372 58812
rect 351920 58760 351972 58812
rect 369124 58760 369176 58812
rect 164608 58692 164660 58744
rect 440240 58692 440292 58744
rect 102232 58624 102284 58676
rect 130568 58624 130620 58676
rect 167000 58624 167052 58676
rect 478880 58624 478932 58676
rect 277952 58556 278004 58608
rect 283564 58556 283616 58608
rect 263416 57196 263468 57248
rect 273260 57196 273312 57248
rect 279424 57196 279476 57248
rect 287060 57196 287112 57248
rect 303160 57196 303212 57248
rect 313188 57196 313240 57248
rect 460204 57196 460256 57248
rect 464896 57196 464948 57248
rect 274732 56924 274784 56976
rect 277768 56924 277820 56976
rect 262220 56516 262272 56568
rect 266360 56516 266412 56568
rect 268844 56516 268896 56568
rect 274272 56516 274324 56568
rect 280988 56516 281040 56568
rect 286324 56516 286376 56568
rect 300308 56516 300360 56568
rect 302240 56516 302292 56568
rect 309784 56516 309836 56568
rect 314292 56516 314344 56568
rect 316684 56516 316736 56568
rect 322204 56516 322256 56568
rect 301320 56448 301372 56500
rect 305920 56448 305972 56500
rect 203524 55836 203576 55888
rect 228364 55836 228416 55888
rect 271144 55836 271196 55888
rect 291844 55836 291896 55888
rect 293960 55836 294012 55888
rect 303528 55836 303580 55888
rect 307668 55836 307720 55888
rect 321468 55836 321520 55888
rect 361672 55836 361724 55888
rect 377404 55836 377456 55888
rect 306104 54748 306156 54800
rect 309876 54748 309928 54800
rect 306012 54680 306064 54732
rect 309784 54680 309836 54732
rect 305736 54612 305788 54664
rect 312544 54612 312596 54664
rect 273260 54544 273312 54596
rect 276112 54544 276164 54596
rect 305644 54544 305696 54596
rect 323768 54544 323820 54596
rect 267004 54476 267056 54528
rect 284300 54476 284352 54528
rect 287060 54476 287112 54528
rect 319444 54476 319496 54528
rect 315396 54340 315448 54392
rect 318340 54340 318392 54392
rect 291936 54136 291988 54188
rect 299112 54136 299164 54188
rect 287704 54068 287756 54120
rect 295340 54068 295392 54120
rect 410524 54068 410576 54120
rect 413928 54068 413980 54120
rect 266360 53184 266412 53236
rect 280804 53184 280856 53236
rect 295984 53184 296036 53236
rect 309968 53184 310020 53236
rect 265624 53116 265676 53168
rect 272524 53116 272576 53168
rect 274088 53116 274140 53168
rect 297364 53116 297416 53168
rect 321468 53116 321520 53168
rect 330484 53116 330536 53168
rect 261484 53048 261536 53100
rect 273904 53048 273956 53100
rect 273996 52980 274048 53032
rect 297456 53048 297508 53100
rect 326344 53048 326396 53100
rect 350540 53048 350592 53100
rect 274272 52912 274324 52964
rect 276020 52912 276072 52964
rect 302240 51960 302292 52012
rect 305000 51960 305052 52012
rect 422944 51824 422996 51876
rect 428464 51824 428516 51876
rect 315304 51756 315356 51808
rect 320732 51756 320784 51808
rect 284300 51688 284352 51740
rect 290832 51688 290884 51740
rect 303528 51688 303580 51740
rect 311164 51688 311216 51740
rect 314292 51688 314344 51740
rect 320824 51688 320876 51740
rect 210424 51620 210476 51672
rect 212540 51620 212592 51672
rect 345756 51348 345808 51400
rect 348424 51348 348476 51400
rect 330484 50804 330536 50856
rect 336096 50804 336148 50856
rect 318156 50736 318208 50788
rect 323676 50736 323728 50788
rect 290464 50532 290516 50584
rect 293224 50532 293276 50584
rect 276020 50396 276072 50448
rect 287612 50396 287664 50448
rect 305828 50396 305880 50448
rect 310428 50396 310480 50448
rect 275284 50328 275336 50380
rect 285680 50328 285732 50380
rect 290556 50328 290608 50380
rect 305644 50328 305696 50380
rect 305920 50328 305972 50380
rect 319536 50328 319588 50380
rect 299112 49784 299164 49836
rect 301504 49784 301556 49836
rect 277768 49648 277820 49700
rect 282920 49648 282972 49700
rect 313188 49648 313240 49700
rect 318156 49648 318208 49700
rect 413928 49648 413980 49700
rect 418160 49648 418212 49700
rect 464896 49648 464948 49700
rect 471244 49648 471296 49700
rect 295340 49240 295392 49292
rect 304264 49240 304316 49292
rect 300216 49172 300268 49224
rect 310612 49172 310664 49224
rect 286416 49104 286468 49156
rect 294604 49104 294656 49156
rect 300124 49104 300176 49156
rect 310520 49104 310572 49156
rect 290832 49036 290884 49088
rect 308496 49036 308548 49088
rect 177212 48968 177264 49020
rect 440332 48968 440384 49020
rect 287612 48220 287664 48272
rect 291936 48220 291988 48272
rect 318064 48220 318116 48272
rect 323584 48220 323636 48272
rect 318340 48152 318392 48204
rect 321008 48152 321060 48204
rect 276664 47676 276716 47728
rect 282184 47676 282236 47728
rect 276112 47608 276164 47660
rect 284944 47608 284996 47660
rect 269764 47540 269816 47592
rect 283656 47540 283708 47592
rect 285680 47540 285732 47592
rect 293868 47540 293920 47592
rect 305000 47540 305052 47592
rect 309600 47540 309652 47592
rect 458824 47540 458876 47592
rect 461308 47540 461360 47592
rect 467196 47540 467248 47592
rect 476764 47540 476816 47592
rect 118424 46860 118476 46912
rect 580172 46860 580224 46912
rect 310520 46792 310572 46844
rect 313280 46792 313332 46844
rect 319444 46792 319496 46844
rect 322848 46792 322900 46844
rect 310612 46724 310664 46776
rect 313464 46724 313516 46776
rect 282920 46180 282972 46232
rect 290648 46180 290700 46232
rect 303068 46180 303120 46232
rect 308404 46180 308456 46232
rect 310428 46180 310480 46232
rect 316776 46180 316828 46232
rect 320732 46180 320784 46232
rect 338764 46180 338816 46232
rect 350540 46180 350592 46232
rect 362224 46180 362276 46232
rect 418160 46180 418212 46232
rect 429108 46180 429160 46232
rect 3424 45500 3476 45552
rect 178224 45500 178276 45552
rect 284944 45500 284996 45552
rect 287612 45500 287664 45552
rect 293868 44956 293920 45008
rect 302240 44956 302292 45008
rect 228364 44888 228416 44940
rect 233884 44888 233936 44940
rect 294604 44888 294656 44940
rect 309048 44888 309100 44940
rect 175280 44820 175332 44872
rect 580264 44820 580316 44872
rect 298744 44684 298796 44736
rect 303804 44684 303856 44736
rect 311164 44548 311216 44600
rect 317328 44548 317380 44600
rect 286324 44412 286376 44464
rect 289728 44412 289780 44464
rect 320824 44276 320876 44328
rect 323032 44276 323084 44328
rect 359464 43732 359516 43784
rect 363604 43732 363656 43784
rect 308496 43528 308548 43580
rect 317052 43528 317104 43580
rect 309968 43460 310020 43512
rect 319444 43460 319496 43512
rect 323768 43460 323820 43512
rect 326068 43460 326120 43512
rect 177948 43392 178000 43444
rect 447140 43392 447192 43444
rect 309876 43324 309928 43376
rect 312268 43324 312320 43376
rect 309784 43188 309836 43240
rect 311900 43188 311952 43240
rect 456064 43052 456116 43104
rect 458548 43052 458600 43104
rect 297456 42848 297508 42900
rect 300768 42848 300820 42900
rect 297364 42780 297416 42832
rect 300124 42780 300176 42832
rect 287612 42372 287664 42424
rect 292028 42372 292080 42424
rect 289084 42100 289136 42152
rect 297640 42100 297692 42152
rect 334624 42100 334676 42152
rect 340144 42100 340196 42152
rect 293224 42032 293276 42084
rect 303712 42032 303764 42084
rect 319536 42032 319588 42084
rect 336188 42032 336240 42084
rect 322204 41556 322256 41608
rect 324964 41556 325016 41608
rect 313924 41352 313976 41404
rect 316684 41352 316736 41404
rect 322848 41352 322900 41404
rect 327724 41352 327776 41404
rect 317328 41284 317380 41336
rect 325056 41284 325108 41336
rect 309048 41216 309100 41268
rect 310704 41216 310756 41268
rect 309600 40740 309652 40792
rect 321100 40740 321152 40792
rect 99380 40672 99432 40724
rect 130476 40672 130528 40724
rect 233884 40672 233936 40724
rect 245660 40672 245712 40724
rect 305644 40672 305696 40724
rect 322940 40672 322992 40724
rect 429108 40672 429160 40724
rect 439504 40672 439556 40724
rect 290648 39992 290700 40044
rect 294604 39992 294656 40044
rect 303712 39992 303764 40044
rect 307024 39992 307076 40044
rect 313464 39992 313516 40044
rect 317236 39992 317288 40044
rect 461308 39992 461360 40044
rect 468484 39992 468536 40044
rect 313280 39924 313332 39976
rect 317328 39924 317380 39976
rect 312268 39856 312320 39908
rect 318524 39856 318576 39908
rect 311900 39788 311952 39840
rect 318432 39788 318484 39840
rect 301504 39380 301556 39432
rect 315304 39380 315356 39432
rect 318156 39380 318208 39432
rect 337936 39380 337988 39432
rect 177856 39312 177908 39364
rect 431960 39312 432012 39364
rect 338764 38428 338816 38480
rect 347136 38428 347188 38480
rect 303804 37884 303856 37936
rect 312636 37884 312688 37936
rect 316776 37884 316828 37936
rect 327080 37884 327132 37936
rect 322940 37612 322992 37664
rect 326160 37612 326212 37664
rect 297640 37204 297692 37256
rect 300492 37204 300544 37256
rect 318432 37204 318484 37256
rect 320824 37204 320876 37256
rect 337936 37204 337988 37256
rect 340788 37204 340840 37256
rect 345664 37204 345716 37256
rect 348516 37204 348568 37256
rect 318524 37136 318576 37188
rect 320916 37136 320968 37188
rect 317052 37068 317104 37120
rect 322756 37068 322808 37120
rect 310704 36932 310756 36984
rect 316776 36932 316828 36984
rect 317328 36796 317380 36848
rect 330484 36796 330536 36848
rect 283748 36728 283800 36780
rect 290372 36728 290424 36780
rect 302976 36728 303028 36780
rect 316868 36728 316920 36780
rect 317236 36728 317288 36780
rect 330576 36728 330628 36780
rect 273904 36660 273956 36712
rect 284944 36660 284996 36712
rect 302240 36660 302292 36712
rect 323768 36660 323820 36712
rect 326068 36660 326120 36712
rect 336004 36660 336056 36712
rect 245660 36592 245712 36644
rect 273996 36592 274048 36644
rect 289728 36592 289780 36644
rect 311164 36592 311216 36644
rect 323032 36592 323084 36644
rect 340696 36592 340748 36644
rect 362224 36592 362276 36644
rect 367744 36592 367796 36644
rect 420184 36592 420236 36644
rect 429844 36592 429896 36644
rect 45560 36524 45612 36576
rect 129372 36524 129424 36576
rect 176384 36524 176436 36576
rect 404360 36524 404412 36576
rect 428464 36524 428516 36576
rect 454868 36524 454920 36576
rect 458548 36524 458600 36576
rect 463884 36524 463936 36576
rect 300768 36048 300820 36100
rect 308496 36048 308548 36100
rect 377404 35300 377456 35352
rect 381544 35300 381596 35352
rect 312544 35164 312596 35216
rect 324320 35164 324372 35216
rect 326160 34892 326212 34944
rect 333244 34892 333296 34944
rect 323676 34416 323728 34468
rect 329196 34416 329248 34468
rect 340788 34416 340840 34468
rect 353944 34416 353996 34468
rect 163872 34348 163924 34400
rect 360200 34348 360252 34400
rect 163504 34280 163556 34332
rect 416780 34280 416832 34332
rect 471244 34280 471296 34332
rect 476120 34280 476172 34332
rect 163320 34212 163372 34264
rect 422300 34212 422352 34264
rect 163412 34144 163464 34196
rect 423680 34144 423732 34196
rect 163228 34076 163280 34128
rect 427820 34076 427872 34128
rect 173164 34008 173216 34060
rect 539692 34008 539744 34060
rect 173256 33940 173308 33992
rect 542360 33940 542412 33992
rect 172980 33872 173032 33924
rect 546500 33872 546552 33924
rect 172888 33804 172940 33856
rect 552020 33804 552072 33856
rect 173072 33736 173124 33788
rect 553400 33736 553452 33788
rect 337384 33124 337436 33176
rect 339960 33124 340012 33176
rect 340144 33056 340196 33108
rect 345940 33056 345992 33108
rect 467104 33056 467156 33108
rect 472348 33056 472400 33108
rect 340696 32988 340748 33040
rect 343640 32988 343692 33040
rect 3424 32784 3476 32836
rect 7656 32784 7708 32836
rect 145288 32648 145340 32700
rect 187700 32648 187752 32700
rect 145196 32580 145248 32632
rect 194600 32580 194652 32632
rect 145380 32512 145432 32564
rect 198740 32512 198792 32564
rect 369124 32512 369176 32564
rect 379520 32512 379572 32564
rect 429844 32512 429896 32564
rect 440884 32512 440936 32564
rect 174452 32444 174504 32496
rect 556252 32444 556304 32496
rect 174360 32376 174412 32428
rect 564532 32376 564584 32428
rect 336188 31832 336240 31884
rect 342904 31832 342956 31884
rect 323584 31696 323636 31748
rect 326344 31696 326396 31748
rect 160468 31560 160520 31612
rect 382280 31560 382332 31612
rect 160560 31492 160612 31544
rect 389180 31492 389232 31544
rect 163044 31424 163096 31476
rect 423772 31424 423824 31476
rect 163136 31356 163188 31408
rect 426440 31356 426492 31408
rect 454868 31356 454920 31408
rect 458824 31356 458876 31408
rect 164516 31288 164568 31340
rect 438860 31288 438912 31340
rect 463884 31288 463936 31340
rect 473360 31288 473412 31340
rect 172520 31220 172572 31272
rect 540980 31220 541032 31272
rect 172612 31152 172664 31204
rect 545120 31152 545172 31204
rect 172704 31084 172756 31136
rect 547972 31084 548024 31136
rect 172796 31016 172848 31068
rect 550640 31016 550692 31068
rect 327080 30948 327132 31000
rect 330668 30948 330720 31000
rect 300492 30268 300544 30320
rect 302240 30268 302292 30320
rect 325056 30268 325108 30320
rect 327908 30268 327960 30320
rect 339960 30268 340012 30320
rect 345020 30268 345072 30320
rect 343640 30200 343692 30252
rect 347044 30200 347096 30252
rect 290372 29656 290424 29708
rect 309784 29656 309836 29708
rect 322756 29656 322808 29708
rect 344468 29656 344520 29708
rect 472348 29656 472400 29708
rect 477500 29656 477552 29708
rect 168748 29588 168800 29640
rect 490012 29588 490064 29640
rect 154028 28908 154080 28960
rect 289820 28908 289872 28960
rect 308496 28908 308548 28960
rect 316592 28908 316644 28960
rect 316868 28908 316920 28960
rect 319628 28908 319680 28960
rect 336096 28908 336148 28960
rect 341064 28908 341116 28960
rect 347136 28908 347188 28960
rect 352564 28908 352616 28960
rect 379520 28908 379572 28960
rect 382924 28908 382976 28960
rect 166632 28840 166684 28892
rect 375380 28840 375432 28892
rect 166540 28772 166592 28824
rect 397460 28772 397512 28824
rect 162032 28704 162084 28756
rect 407120 28704 407172 28756
rect 162952 28636 163004 28688
rect 415492 28636 415544 28688
rect 166172 28568 166224 28620
rect 449900 28568 449952 28620
rect 165988 28500 166040 28552
rect 452660 28500 452712 28552
rect 166080 28432 166132 28484
rect 456892 28432 456944 28484
rect 166264 28364 166316 28416
rect 459560 28364 459612 28416
rect 171692 28296 171744 28348
rect 521660 28296 521712 28348
rect 171600 28228 171652 28280
rect 524420 28228 524472 28280
rect 146944 28160 146996 28212
rect 209780 28160 209832 28212
rect 316592 28160 316644 28212
rect 318064 28160 318116 28212
rect 345940 28160 345992 28212
rect 353300 28160 353352 28212
rect 146852 28092 146904 28144
rect 205640 28092 205692 28144
rect 146760 28024 146812 28076
rect 201500 28024 201552 28076
rect 324964 27616 325016 27668
rect 327080 27616 327132 27668
rect 307024 27548 307076 27600
rect 312176 27548 312228 27600
rect 348516 27548 348568 27600
rect 352656 27548 352708 27600
rect 312636 27004 312688 27056
rect 320088 27004 320140 27056
rect 323768 27004 323820 27056
rect 329104 27004 329156 27056
rect 145104 26936 145156 26988
rect 193312 26936 193364 26988
rect 300124 26936 300176 26988
rect 321192 26936 321244 26988
rect 324320 26936 324372 26988
rect 334624 26936 334676 26988
rect 160376 26868 160428 26920
rect 385040 26868 385092 26920
rect 439504 26868 439556 26920
rect 446404 26868 446456 26920
rect 464344 26868 464396 26920
rect 493324 26868 493376 26920
rect 302240 26324 302292 26376
rect 306380 26324 306432 26376
rect 283564 26120 283616 26172
rect 292764 26120 292816 26172
rect 145012 26052 145064 26104
rect 186320 26052 186372 26104
rect 283656 26052 283708 26104
rect 294052 26052 294104 26104
rect 363604 26052 363656 26104
rect 367560 26052 367612 26104
rect 152740 25984 152792 26036
rect 253940 25984 253992 26036
rect 280804 25984 280856 26036
rect 294144 25984 294196 26036
rect 315304 25984 315356 26036
rect 320180 25984 320232 26036
rect 321100 25984 321152 26036
rect 329012 25984 329064 26036
rect 333244 25984 333296 26036
rect 343640 25984 343692 26036
rect 349804 25984 349856 26036
rect 364984 25984 365036 26036
rect 162584 25916 162636 25968
rect 368480 25916 368532 25968
rect 162492 25848 162544 25900
rect 390560 25848 390612 25900
rect 170220 25780 170272 25832
rect 506480 25780 506532 25832
rect 171508 25712 171560 25764
rect 528560 25712 528612 25764
rect 174176 25644 174228 25696
rect 558920 25644 558972 25696
rect 174084 25576 174136 25628
rect 563060 25576 563112 25628
rect 174268 25508 174320 25560
rect 565820 25508 565872 25560
rect 302884 24828 302936 24880
rect 307116 24828 307168 24880
rect 321008 24828 321060 24880
rect 323584 24828 323636 24880
rect 291844 24556 291896 24608
rect 294328 24556 294380 24608
rect 316776 24420 316828 24472
rect 319536 24420 319588 24472
rect 440884 24284 440936 24336
rect 443736 24284 443788 24336
rect 292028 24216 292080 24268
rect 300676 24216 300728 24268
rect 273996 24148 274048 24200
rect 292672 24148 292724 24200
rect 320088 24148 320140 24200
rect 324964 24148 325016 24200
rect 327908 24148 327960 24200
rect 344376 24148 344428 24200
rect 2964 24080 3016 24132
rect 189172 24080 189224 24132
rect 284944 24080 284996 24132
rect 304448 24080 304500 24132
rect 326344 24080 326396 24132
rect 342260 24080 342312 24132
rect 344468 24080 344520 24132
rect 349896 24080 349948 24132
rect 353300 24080 353352 24132
rect 359280 24080 359332 24132
rect 141240 23400 141292 23452
rect 142160 23400 142212 23452
rect 146668 23400 146720 23452
rect 204260 23400 204312 23452
rect 381544 23400 381596 23452
rect 384304 23400 384356 23452
rect 146484 23332 146536 23384
rect 208400 23332 208452 23384
rect 146576 23264 146628 23316
rect 211160 23264 211212 23316
rect 272524 23264 272576 23316
rect 275008 23264 275060 23316
rect 309784 23264 309836 23316
rect 312912 23264 312964 23316
rect 152464 23196 152516 23248
rect 273260 23196 273312 23248
rect 308404 23196 308456 23248
rect 313280 23196 313332 23248
rect 152372 23128 152424 23180
rect 280160 23128 280212 23180
rect 142620 23060 142672 23112
rect 149060 23060 149112 23112
rect 153752 23060 153804 23112
rect 291200 23060 291252 23112
rect 141332 22992 141384 23044
rect 145012 22992 145064 23044
rect 153936 22992 153988 23044
rect 293960 22992 294012 23044
rect 294604 22992 294656 23044
rect 305644 22992 305696 23044
rect 153844 22924 153896 22976
rect 300860 22924 300912 22976
rect 3424 22856 3476 22908
rect 178132 22856 178184 22908
rect 291936 22856 291988 22908
rect 307024 22856 307076 22908
rect 129648 22788 129700 22840
rect 305000 22788 305052 22840
rect 306380 22788 306432 22840
rect 340052 22788 340104 22840
rect 341064 22788 341116 22840
rect 358084 22788 358136 22840
rect 120724 22720 120776 22772
rect 580264 22720 580316 22772
rect 329012 22652 329064 22704
rect 334808 22652 334860 22704
rect 312176 22312 312228 22364
rect 315304 22312 315356 22364
rect 294328 22040 294380 22092
rect 298008 22040 298060 22092
rect 352656 22040 352708 22092
rect 357164 22040 357216 22092
rect 446404 22040 446456 22092
rect 448888 22040 448940 22092
rect 329196 21700 329248 21752
rect 341524 21700 341576 21752
rect 327080 21632 327132 21684
rect 340144 21632 340196 21684
rect 344284 21632 344336 21684
rect 352656 21632 352708 21684
rect 177672 21564 177724 21616
rect 418160 21564 418212 21616
rect 169944 21496 169996 21548
rect 506572 21496 506624 21548
rect 170128 21428 170180 21480
rect 509240 21428 509292 21480
rect 170036 21360 170088 21412
rect 513380 21360 513432 21412
rect 150900 20612 150952 20664
rect 255320 20612 255372 20664
rect 300676 20612 300728 20664
rect 308496 20612 308548 20664
rect 347044 20612 347096 20664
rect 349804 20612 349856 20664
rect 349896 20612 349948 20664
rect 355600 20612 355652 20664
rect 359280 20612 359332 20664
rect 365076 20612 365128 20664
rect 367560 20612 367612 20664
rect 371240 20612 371292 20664
rect 526444 20612 526496 20664
rect 579988 20612 580040 20664
rect 150992 20544 151044 20596
rect 259552 20544 259604 20596
rect 151084 20476 151136 20528
rect 262220 20476 262272 20528
rect 151176 20408 151228 20460
rect 269120 20408 269172 20460
rect 275008 20408 275060 20460
rect 288348 20408 288400 20460
rect 292672 20408 292724 20460
rect 300124 20408 300176 20460
rect 152280 20340 152332 20392
rect 276020 20340 276072 20392
rect 292764 20340 292816 20392
rect 307208 20340 307260 20392
rect 153660 20272 153712 20324
rect 298100 20272 298152 20324
rect 312912 20272 312964 20324
rect 327080 20272 327132 20324
rect 161940 20204 161992 20256
rect 402980 20204 403032 20256
rect 170956 20136 171008 20188
rect 488540 20136 488592 20188
rect 168656 20068 168708 20120
rect 495440 20068 495492 20120
rect 168564 20000 168616 20052
rect 498292 20000 498344 20052
rect 120080 19932 120132 19984
rect 139676 19932 139728 19984
rect 171416 19932 171468 19984
rect 531412 19932 531464 19984
rect 149704 19864 149756 19916
rect 237380 19864 237432 19916
rect 330668 19252 330720 19304
rect 334716 19252 334768 19304
rect 330576 18776 330628 18828
rect 338764 18776 338816 18828
rect 448888 18776 448940 18828
rect 452752 18776 452804 18828
rect 294052 18708 294104 18760
rect 304356 18708 304408 18760
rect 146208 18640 146260 18692
rect 218060 18640 218112 18692
rect 298008 18640 298060 18692
rect 312544 18640 312596 18692
rect 330484 18640 330536 18692
rect 339316 18640 339368 18692
rect 340144 18640 340196 18692
rect 349160 18640 349212 18692
rect 357164 18640 357216 18692
rect 369124 18640 369176 18692
rect 173992 18572 174044 18624
rect 560300 18572 560352 18624
rect 443736 17892 443788 17944
rect 449164 17892 449216 17944
rect 288348 17688 288400 17740
rect 297364 17688 297416 17740
rect 148232 17620 148284 17672
rect 226340 17620 226392 17672
rect 294144 17620 294196 17672
rect 312636 17620 312688 17672
rect 355600 17620 355652 17672
rect 365720 17620 365772 17672
rect 367744 17620 367796 17672
rect 377404 17620 377456 17672
rect 161848 17552 161900 17604
rect 398932 17552 398984 17604
rect 164424 17484 164476 17536
rect 436100 17484 436152 17536
rect 164332 17416 164384 17468
rect 441620 17416 441672 17468
rect 165896 17348 165948 17400
rect 462320 17348 462372 17400
rect 171324 17280 171376 17332
rect 523040 17280 523092 17332
rect 171232 17212 171284 17264
rect 527180 17212 527232 17264
rect 342260 16804 342312 16856
rect 346400 16804 346452 16856
rect 304448 16260 304500 16312
rect 308404 16260 308456 16312
rect 149612 15920 149664 15972
rect 248420 15920 248472 15972
rect 323584 15920 323636 15972
rect 333244 15920 333296 15972
rect 334808 15920 334860 15972
rect 339040 15920 339092 15972
rect 342904 15920 342956 15972
rect 347872 15920 347924 15972
rect 35992 15852 36044 15904
rect 124864 15852 124916 15904
rect 176292 15852 176344 15904
rect 411904 15852 411956 15904
rect 349804 15716 349856 15768
rect 352288 15716 352340 15768
rect 452752 15580 452804 15632
rect 458180 15580 458232 15632
rect 152096 15104 152148 15156
rect 276112 15104 276164 15156
rect 152188 15036 152240 15088
rect 279056 15036 279108 15088
rect 308496 15036 308548 15088
rect 319812 15036 319864 15088
rect 339316 15036 339368 15088
rect 342812 15036 342864 15088
rect 152004 14968 152056 15020
rect 283104 14968 283156 15020
rect 300124 14968 300176 15020
rect 314752 14968 314804 15020
rect 334624 14968 334676 15020
rect 340236 14968 340288 15020
rect 365076 14968 365128 15020
rect 370504 14968 370556 15020
rect 153568 14900 153620 14952
rect 297272 14900 297324 14952
rect 304264 14900 304316 14952
rect 320732 14900 320784 14952
rect 324964 14900 325016 14952
rect 347136 14900 347188 14952
rect 160100 14832 160152 14884
rect 384304 14832 384356 14884
rect 160192 14764 160244 14816
rect 387800 14764 387852 14816
rect 160284 14696 160336 14748
rect 390652 14696 390704 14748
rect 161756 14628 161808 14680
rect 400864 14628 400916 14680
rect 162860 14560 162912 14612
rect 420920 14560 420972 14612
rect 449164 14560 449216 14612
rect 454592 14560 454644 14612
rect 165804 14492 165856 14544
rect 459192 14492 459244 14544
rect 468484 14492 468536 14544
rect 482284 14492 482336 14544
rect 174820 14424 174872 14476
rect 567568 14424 567620 14476
rect 150808 14356 150860 14408
rect 264980 14356 265032 14408
rect 348424 14356 348476 14408
rect 350908 14356 350960 14408
rect 150716 14288 150768 14340
rect 261760 14288 261812 14340
rect 147036 14220 147088 14272
rect 190460 14220 190512 14272
rect 364984 13880 365036 13932
rect 367744 13880 367796 13932
rect 319444 13812 319496 13864
rect 322204 13812 322256 13864
rect 321192 13744 321244 13796
rect 326344 13744 326396 13796
rect 353944 13744 353996 13796
rect 356704 13744 356756 13796
rect 479524 13744 479576 13796
rect 481732 13744 481784 13796
rect 341524 13676 341576 13728
rect 347044 13676 347096 13728
rect 329104 13200 329156 13252
rect 334624 13200 334676 13252
rect 493324 13064 493376 13116
rect 507860 13064 507912 13116
rect 340052 12452 340104 12504
rect 342996 12452 343048 12504
rect 146392 12384 146444 12436
rect 214472 12384 214524 12436
rect 358084 12384 358136 12436
rect 361580 12384 361632 12436
rect 458824 12384 458876 12436
rect 461676 12384 461728 12436
rect 148140 12316 148192 12368
rect 222752 12316 222804 12368
rect 147956 12248 148008 12300
rect 226432 12248 226484 12300
rect 307116 12248 307168 12300
rect 311900 12248 311952 12300
rect 148048 12180 148100 12232
rect 229376 12180 229428 12232
rect 149520 12112 149572 12164
rect 240140 12112 240192 12164
rect 320732 12112 320784 12164
rect 149428 12044 149480 12096
rect 242900 12044 242952 12096
rect 319628 12044 319680 12096
rect 322296 12044 322348 12096
rect 352656 12112 352708 12164
rect 357532 12112 357584 12164
rect 329104 12044 329156 12096
rect 347872 12044 347924 12096
rect 359464 12044 359516 12096
rect 165160 11976 165212 12028
rect 382372 11976 382424 12028
rect 382924 11976 382976 12028
rect 389824 11976 389876 12028
rect 161664 11908 161716 11960
rect 402520 11908 402572 11960
rect 161572 11840 161624 11892
rect 406016 11840 406068 11892
rect 165712 11772 165764 11824
rect 455696 11772 455748 11824
rect 476764 11772 476816 11824
rect 479524 11772 479576 11824
rect 126980 11704 127032 11756
rect 128176 11704 128228 11756
rect 135260 11704 135312 11756
rect 136456 11704 136508 11756
rect 169852 11704 169904 11756
rect 511264 11704 511316 11756
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 226340 11636 226392 11688
rect 227536 11636 227588 11688
rect 259460 11636 259512 11688
rect 260656 11636 260708 11688
rect 311164 11636 311216 11688
rect 314660 11636 314712 11688
rect 327724 11636 327776 11688
rect 330484 11636 330536 11688
rect 316684 10956 316736 11008
rect 319444 10956 319496 11008
rect 339040 10956 339092 11008
rect 342720 10956 342772 11008
rect 347136 10956 347188 11008
rect 349252 10956 349304 11008
rect 318064 10888 318116 10940
rect 322388 10888 322440 10940
rect 112352 10684 112404 10736
rect 138388 10684 138440 10736
rect 92480 10616 92532 10668
rect 130384 10616 130436 10668
rect 89168 10548 89220 10600
rect 137008 10548 137060 10600
rect 75000 10480 75052 10532
rect 134524 10480 134576 10532
rect 71504 10412 71556 10464
rect 135904 10412 135956 10464
rect 20168 10344 20220 10396
rect 95884 10344 95936 10396
rect 106464 10344 106516 10396
rect 138480 10344 138532 10396
rect 350908 10344 350960 10396
rect 363512 10344 363564 10396
rect 365720 10344 365772 10396
rect 374092 10344 374144 10396
rect 458180 10344 458232 10396
rect 465724 10344 465776 10396
rect 56784 10276 56836 10328
rect 134340 10276 134392 10328
rect 169760 10276 169812 10328
rect 503720 10276 503772 10328
rect 307208 9596 307260 9648
rect 309324 9596 309376 9648
rect 320916 9596 320968 9648
rect 324688 9596 324740 9648
rect 336004 9596 336056 9648
rect 342168 9596 342220 9648
rect 320824 9528 320876 9580
rect 324780 9528 324832 9580
rect 109316 9392 109368 9444
rect 138296 9392 138348 9444
rect 82084 9324 82136 9376
rect 136916 9324 136968 9376
rect 77392 9256 77444 9308
rect 135720 9256 135772 9308
rect 73804 9188 73856 9240
rect 135628 9188 135680 9240
rect 177488 9188 177540 9240
rect 207388 9188 207440 9240
rect 70308 9120 70360 9172
rect 135812 9120 135864 9172
rect 146300 9120 146352 9172
rect 210976 9120 211028 9172
rect 352288 9120 352340 9172
rect 364616 9120 364668 9172
rect 43076 9052 43128 9104
rect 122104 9052 122156 9104
rect 149336 9052 149388 9104
rect 247592 9052 247644 9104
rect 282184 9052 282236 9104
rect 302148 9052 302200 9104
rect 304356 9052 304408 9104
rect 312268 9052 312320 9104
rect 315304 9052 315356 9104
rect 330760 9052 330812 9104
rect 338764 9052 338816 9104
rect 351460 9052 351512 9104
rect 361580 9052 361632 9104
rect 377680 9052 377732 9104
rect 53748 8984 53800 9036
rect 134248 8984 134300 9036
rect 161480 8984 161532 9036
rect 407212 8984 407264 9036
rect 14740 8916 14792 8968
rect 131764 8916 131816 8968
rect 168472 8916 168524 8968
rect 493508 8916 493560 8968
rect 507860 8916 507912 8968
rect 526628 8916 526680 8968
rect 312636 8304 312688 8356
rect 316224 8304 316276 8356
rect 297364 8236 297416 8288
rect 303528 8236 303580 8288
rect 377404 8236 377456 8288
rect 379980 8236 380032 8288
rect 135260 8100 135312 8152
rect 135444 8100 135496 8152
rect 123484 7896 123536 7948
rect 139584 7896 139636 7948
rect 66720 7828 66772 7880
rect 135536 7828 135588 7880
rect 52552 7760 52604 7812
rect 134064 7760 134116 7812
rect 50160 7692 50212 7744
rect 134156 7692 134208 7744
rect 312544 7692 312596 7744
rect 323308 7692 323360 7744
rect 28908 7624 28960 7676
rect 126336 7624 126388 7676
rect 314752 7624 314804 7676
rect 327080 7624 327132 7676
rect 334716 7624 334768 7676
rect 356336 7624 356388 7676
rect 15936 7556 15988 7608
rect 131672 7556 131724 7608
rect 164240 7556 164292 7608
rect 443828 7556 443880 7608
rect 454592 7556 454644 7608
rect 473452 7556 473504 7608
rect 311900 7488 311952 7540
rect 317420 7488 317472 7540
rect 149980 6808 150032 6860
rect 203892 6808 203944 6860
rect 149244 6740 149296 6792
rect 246396 6740 246448 6792
rect 150624 6672 150676 6724
rect 267740 6672 267792 6724
rect 151820 6604 151872 6656
rect 278320 6604 278372 6656
rect 40684 6536 40736 6588
rect 132684 6536 132736 6588
rect 151912 6536 151964 6588
rect 281908 6536 281960 6588
rect 333244 6536 333296 6588
rect 338672 6536 338724 6588
rect 38384 6468 38436 6520
rect 133052 6468 133104 6520
rect 153476 6468 153528 6520
rect 292580 6468 292632 6520
rect 324688 6468 324740 6520
rect 334072 6468 334124 6520
rect 37188 6400 37240 6452
rect 132776 6400 132828 6452
rect 153384 6400 153436 6452
rect 296076 6400 296128 6452
rect 324780 6400 324832 6452
rect 333980 6400 334032 6452
rect 340236 6400 340288 6452
rect 352840 6400 352892 6452
rect 33600 6332 33652 6384
rect 132960 6332 133012 6384
rect 153292 6332 153344 6384
rect 299664 6332 299716 6384
rect 330760 6332 330812 6384
rect 343640 6332 343692 6384
rect 31300 6264 31352 6316
rect 133144 6264 133196 6316
rect 153200 6264 153252 6316
rect 300768 6264 300820 6316
rect 305644 6264 305696 6316
rect 309232 6264 309284 6316
rect 309324 6264 309376 6316
rect 339868 6264 339920 6316
rect 342996 6264 343048 6316
rect 357164 6264 357216 6316
rect 30104 6196 30156 6248
rect 132868 6196 132920 6248
rect 175188 6196 175240 6248
rect 573916 6196 573968 6248
rect 24216 6128 24268 6180
rect 131580 6128 131632 6180
rect 176568 6128 176620 6180
rect 578608 6128 578660 6180
rect 144920 6060 144972 6112
rect 196808 6060 196860 6112
rect 356704 5924 356756 5976
rect 362960 5924 363012 5976
rect 351460 5856 351512 5908
rect 353300 5856 353352 5908
rect 319536 5516 319588 5568
rect 324412 5516 324464 5568
rect 326344 5516 326396 5568
rect 332692 5516 332744 5568
rect 479524 5516 479576 5568
rect 482836 5516 482888 5568
rect 143816 5380 143868 5432
rect 149244 5380 149296 5432
rect 122288 5312 122340 5364
rect 139952 5312 140004 5364
rect 110512 5244 110564 5296
rect 129188 5244 129240 5296
rect 108120 5176 108172 5228
rect 138204 5176 138256 5228
rect 142344 5176 142396 5228
rect 155408 5176 155460 5228
rect 104532 5108 104584 5160
rect 138940 5108 138992 5160
rect 142436 5108 142488 5160
rect 157800 5108 157852 5160
rect 56048 5040 56100 5092
rect 134432 5040 134484 5092
rect 143908 5040 143960 5092
rect 169576 5040 169628 5092
rect 23020 4972 23072 5024
rect 131396 4972 131448 5024
rect 144000 4972 144052 5024
rect 173164 4972 173216 5024
rect 19432 4904 19484 4956
rect 129280 4904 129332 4956
rect 147864 4904 147916 4956
rect 220452 4972 220504 5024
rect 21824 4836 21876 4888
rect 131304 4836 131356 4888
rect 142528 4836 142580 4888
rect 158904 4836 158956 4888
rect 169668 4836 169720 4888
rect 494704 4836 494756 4888
rect 18236 4768 18288 4820
rect 131488 4768 131540 4820
rect 144092 4768 144144 4820
rect 170772 4768 170824 4820
rect 171140 4768 171192 4820
rect 533712 4768 533764 4820
rect 6460 4088 6512 4140
rect 7564 4088 7616 4140
rect 140964 4088 141016 4140
rect 144736 4088 144788 4140
rect 148416 4088 148468 4140
rect 153016 4088 153068 4140
rect 125876 4020 125928 4072
rect 139768 4020 139820 4072
rect 147772 4020 147824 4072
rect 225144 4088 225196 4140
rect 343640 4088 343692 4140
rect 351644 4088 351696 4140
rect 352564 4088 352616 4140
rect 355232 4088 355284 4140
rect 357164 4088 357216 4140
rect 367008 4088 367060 4140
rect 389824 4088 389876 4140
rect 394240 4088 394292 4140
rect 156696 4020 156748 4072
rect 228732 4020 228784 4072
rect 303528 4020 303580 4072
rect 310244 4020 310296 4072
rect 344376 4020 344428 4072
rect 358728 4020 358780 4072
rect 86868 3952 86920 4004
rect 137284 3952 137336 4004
rect 149152 3952 149204 4004
rect 239312 3952 239364 4004
rect 251180 3952 251232 4004
rect 252376 3952 252428 4004
rect 307024 3952 307076 4004
rect 318524 3952 318576 4004
rect 322388 3952 322440 4004
rect 329196 3952 329248 4004
rect 353300 3952 353352 4004
rect 374000 4020 374052 4072
rect 69112 3884 69164 3936
rect 135352 3884 135404 3936
rect 150440 3884 150492 3936
rect 258264 3884 258316 3936
rect 276020 3884 276072 3936
rect 276756 3884 276808 3936
rect 317420 3884 317472 3936
rect 330392 3884 330444 3936
rect 333980 3884 334032 3936
rect 340972 3884 341024 3936
rect 342812 3884 342864 3936
rect 370228 3952 370280 4004
rect 370504 3952 370556 4004
rect 378876 3952 378928 4004
rect 369124 3884 369176 3936
rect 372896 3884 372948 3936
rect 62028 3816 62080 3868
rect 129004 3816 129056 3868
rect 144460 3816 144512 3868
rect 160100 3816 160152 3868
rect 166724 3816 166776 3868
rect 458088 3816 458140 3868
rect 461676 3816 461728 3868
rect 471060 3816 471112 3868
rect 9956 3748 10008 3800
rect 88892 3748 88944 3800
rect 93952 3748 94004 3800
rect 137100 3748 137152 3800
rect 143448 3748 143500 3800
rect 151820 3748 151872 3800
rect 176108 3748 176160 3800
rect 472256 3748 472308 3800
rect 39580 3680 39632 3732
rect 129096 3680 129148 3732
rect 140688 3680 140740 3732
rect 161296 3680 161348 3732
rect 177580 3680 177632 3732
rect 480536 3680 480588 3732
rect 17040 3612 17092 3664
rect 131948 3612 132000 3664
rect 143724 3612 143776 3664
rect 167184 3612 167236 3664
rect 177396 3612 177448 3664
rect 181444 3612 181496 3664
rect 185584 3612 185636 3664
rect 487620 3612 487672 3664
rect 1676 3544 1728 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 5264 3544 5316 3596
rect 10324 3544 10376 3596
rect 11060 3544 11112 3596
rect 11980 3544 12032 3596
rect 13544 3544 13596 3596
rect 131212 3544 131264 3596
rect 141056 3544 141108 3596
rect 147128 3544 147180 3596
rect 149244 3544 149296 3596
rect 174268 3544 174320 3596
rect 177304 3544 177356 3596
rect 491116 3544 491168 3596
rect 126244 3476 126296 3528
rect 131764 3476 131816 3528
rect 140044 3476 140096 3528
rect 143632 3476 143684 3528
rect 171968 3476 172020 3528
rect 176200 3476 176252 3528
rect 177856 3476 177908 3528
rect 177948 3476 178000 3528
rect 505376 3476 505428 3528
rect 506480 3476 506532 3528
rect 507308 3476 507360 3528
rect 531320 3476 531372 3528
rect 532148 3476 532200 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 572 3408 624 3460
rect 127624 3408 127676 3460
rect 132960 3408 133012 3460
rect 140136 3408 140188 3460
rect 144552 3408 144604 3460
rect 175464 3408 175516 3460
rect 177764 3408 177816 3460
rect 508872 3408 508924 3460
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 147680 3340 147732 3392
rect 156696 3340 156748 3392
rect 141516 3272 141568 3324
rect 143540 3272 143592 3324
rect 147220 3204 147272 3256
rect 189724 3340 189776 3392
rect 218060 3340 218112 3392
rect 219256 3340 219308 3392
rect 242900 3340 242952 3392
rect 244096 3340 244148 3392
rect 302148 3340 302200 3392
rect 309048 3340 309100 3392
rect 322296 3340 322348 3392
rect 325608 3340 325660 3392
rect 329104 3340 329156 3392
rect 336280 3340 336332 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 374092 3340 374144 3392
rect 375288 3340 375340 3392
rect 382372 3340 382424 3392
rect 383568 3340 383620 3392
rect 390652 3340 390704 3392
rect 391848 3340 391900 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 431960 3340 432012 3392
rect 433248 3340 433300 3392
rect 465724 3340 465776 3392
rect 469864 3340 469916 3392
rect 175924 3272 175976 3324
rect 177948 3272 178000 3324
rect 171876 3204 171928 3256
rect 176660 3204 176712 3256
rect 142252 3136 142304 3188
rect 150624 3136 150676 3188
rect 172060 3068 172112 3120
rect 186136 3272 186188 3324
rect 319812 3272 319864 3324
rect 322112 3272 322164 3324
rect 334072 3272 334124 3324
rect 337476 3272 337528 3324
rect 322204 3204 322256 3256
rect 326804 3204 326856 3256
rect 384396 3204 384448 3256
rect 387156 3204 387208 3256
rect 309232 3136 309284 3188
rect 317328 3136 317380 3188
rect 482284 3136 482336 3188
rect 485228 3136 485280 3188
rect 327080 3068 327132 3120
rect 331588 3068 331640 3120
rect 347044 3068 347096 3120
rect 354036 3068 354088 3120
rect 140044 3000 140096 3052
rect 141148 3000 141200 3052
rect 145564 3000 145616 3052
rect 154212 3000 154264 3052
rect 175556 3000 175608 3052
rect 185584 3000 185636 3052
rect 330484 3000 330536 3052
rect 333888 3000 333940 3052
rect 362960 3000 363012 3052
rect 365812 3000 365864 3052
rect 308404 2932 308456 2984
rect 311440 2932 311492 2984
rect 407120 1776 407172 1828
rect 408408 1776 408460 1828
rect 415400 1776 415452 1828
rect 416688 1776 416740 1828
rect 440240 1776 440292 1828
rect 441528 1776 441580 1828
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 527912 3386 527921
rect 3330 527847 3332 527856
rect 3384 527847 3386 527856
rect 3332 527818 3384 527824
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 3068 462398 3096 462567
rect 3056 462392 3108 462398
rect 3056 462334 3108 462340
rect 2962 449576 3018 449585
rect 2962 449511 3018 449520
rect 2976 448594 3004 449511
rect 2964 448588 3016 448594
rect 2964 448530 3016 448536
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3344 422346 3372 423535
rect 3332 422340 3384 422346
rect 3332 422282 3384 422288
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3146 319288 3202 319297
rect 3146 319223 3202 319232
rect 3160 318850 3188 319223
rect 3148 318844 3200 318850
rect 3148 318786 3200 318792
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3344 305046 3372 306167
rect 3332 305040 3384 305046
rect 3332 304982 3384 304988
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3252 266422 3280 267135
rect 3240 266416 3292 266422
rect 3240 266358 3292 266364
rect 2870 254144 2926 254153
rect 2870 254079 2926 254088
rect 2884 253978 2912 254079
rect 2872 253972 2924 253978
rect 2872 253914 2924 253920
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3344 201550 3372 201855
rect 3332 201544 3384 201550
rect 3332 201486 3384 201492
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3344 187746 3372 188799
rect 3332 187740 3384 187746
rect 3332 187682 3384 187688
rect 3332 162920 3384 162926
rect 3330 162888 3332 162897
rect 3384 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3344 84250 3372 84623
rect 3332 84244 3384 84250
rect 3332 84186 3384 84192
rect 3436 79257 3464 606047
rect 3528 149938 3556 671191
rect 3606 619168 3662 619177
rect 3606 619103 3662 619112
rect 3516 149932 3568 149938
rect 3516 149874 3568 149880
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3528 148374 3556 149767
rect 3516 148368 3568 148374
rect 3516 148310 3568 148316
rect 3620 146946 3648 619103
rect 3790 566944 3846 566953
rect 3790 566879 3846 566888
rect 3698 501800 3754 501809
rect 3698 501735 3754 501744
rect 3608 146940 3660 146946
rect 3608 146882 3660 146888
rect 3608 139460 3660 139466
rect 3608 139402 3660 139408
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3528 136678 3556 136711
rect 3516 136672 3568 136678
rect 3516 136614 3568 136620
rect 3620 122834 3648 139402
rect 3528 122806 3648 122834
rect 3528 97617 3556 122806
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3712 80034 3740 501735
rect 3804 160750 3832 566879
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3896 461650 3924 475623
rect 3884 461644 3936 461650
rect 3884 461586 3936 461592
rect 3882 358456 3938 358465
rect 3882 358391 3938 358400
rect 3792 160744 3844 160750
rect 3792 160686 3844 160692
rect 3792 149932 3844 149938
rect 3792 149874 3844 149880
rect 3804 145586 3832 149874
rect 3792 145580 3844 145586
rect 3792 145522 3844 145528
rect 3896 142934 3924 358391
rect 3974 293176 4030 293185
rect 3974 293111 4030 293120
rect 3884 142928 3936 142934
rect 3884 142870 3936 142876
rect 3700 80028 3752 80034
rect 3700 79970 3752 79976
rect 3988 79354 4016 293111
rect 4066 241088 4122 241097
rect 4066 241023 4122 241032
rect 4080 84194 4108 241023
rect 4816 118658 4844 683674
rect 4804 118652 4856 118658
rect 4804 118594 4856 118600
rect 4080 84166 4200 84194
rect 4172 84130 4200 84166
rect 4080 84102 4200 84130
rect 3976 79348 4028 79354
rect 3976 79290 4028 79296
rect 3422 79248 3478 79257
rect 3422 79183 3478 79192
rect 4080 78577 4108 84102
rect 6932 79665 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 7564 632120 7616 632126
rect 7564 632062 7616 632068
rect 7576 120086 7604 632062
rect 17224 579692 17276 579698
rect 17224 579634 17276 579640
rect 8944 527876 8996 527882
rect 8944 527818 8996 527824
rect 7656 136740 7708 136746
rect 7656 136682 7708 136688
rect 7564 120080 7616 120086
rect 7564 120022 7616 120028
rect 6918 79656 6974 79665
rect 6918 79591 6974 79600
rect 4066 78568 4122 78577
rect 4066 78503 4122 78512
rect 6918 75168 6974 75177
rect 6918 75103 6974 75112
rect 3424 71664 3476 71670
rect 3422 71632 3424 71641
rect 3476 71632 3478 71641
rect 3422 71567 3478 71576
rect 3424 69896 3476 69902
rect 3424 69838 3476 69844
rect 2780 69692 2832 69698
rect 2780 69634 2832 69640
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3538
rect 2792 3534 2820 69634
rect 2872 66904 2924 66910
rect 2872 66846 2924 66852
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 66846
rect 3436 58585 3464 69838
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 32836 3476 32842
rect 3424 32778 3476 32784
rect 3436 32473 3464 32778
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 2964 24132 3016 24138
rect 2964 24074 3016 24080
rect 2976 19417 3004 24074
rect 3424 22908 3476 22914
rect 3424 22850 3476 22856
rect 2962 19408 3018 19417
rect 2962 19343 3018 19352
rect 3436 6497 3464 22850
rect 6932 16574 6960 75103
rect 7564 61396 7616 61402
rect 7564 61338 7616 61344
rect 6932 16546 7512 16574
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5276 480 5304 3538
rect 6472 480 6500 4082
rect 7484 3482 7512 16546
rect 7576 4146 7604 61338
rect 7668 32842 7696 136682
rect 8956 122806 8984 527818
rect 10324 422340 10376 422346
rect 10324 422282 10376 422288
rect 9036 135312 9088 135318
rect 9036 135254 9088 135260
rect 8944 122800 8996 122806
rect 8944 122742 8996 122748
rect 8298 72448 8354 72457
rect 8298 72383 8354 72392
rect 7656 32836 7708 32842
rect 7656 32778 7708 32784
rect 8312 16574 8340 72383
rect 9048 71670 9076 135254
rect 10336 126954 10364 422282
rect 13084 318844 13136 318850
rect 13084 318786 13136 318792
rect 13096 129742 13124 318786
rect 14464 162920 14516 162926
rect 14464 162862 14516 162868
rect 14476 133890 14504 162862
rect 14464 133884 14516 133890
rect 14464 133826 14516 133832
rect 13084 129736 13136 129742
rect 13084 129678 13136 129684
rect 10324 126948 10376 126954
rect 10324 126890 10376 126896
rect 17236 121446 17264 579634
rect 18604 266416 18656 266422
rect 18604 266358 18656 266364
rect 18616 131102 18644 266358
rect 23492 144294 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 31024 213988 31076 213994
rect 31024 213930 31076 213936
rect 23480 144288 23532 144294
rect 23480 144230 23532 144236
rect 21364 133952 21416 133958
rect 21364 133894 21416 133900
rect 18604 131096 18656 131102
rect 18604 131038 18656 131044
rect 17224 121440 17276 121446
rect 17224 121382 17276 121388
rect 21376 111790 21404 133894
rect 31036 132462 31064 213930
rect 31024 132456 31076 132462
rect 31024 132398 31076 132404
rect 40052 117298 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 48964 461644 49016 461650
rect 48964 461586 49016 461592
rect 48976 124166 49004 461586
rect 48964 124160 49016 124166
rect 48964 124102 49016 124108
rect 40040 117292 40092 117298
rect 40040 117234 40092 117240
rect 21364 111784 21416 111790
rect 21364 111726 21416 111732
rect 71792 79529 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 84844 448588 84896 448594
rect 84844 448530 84896 448536
rect 71778 79520 71834 79529
rect 71778 79455 71834 79464
rect 84856 78946 84884 448530
rect 84936 371272 84988 371278
rect 84936 371214 84988 371220
rect 84948 128314 84976 371214
rect 88352 141506 88380 702406
rect 105464 699718 105492 703520
rect 137848 700330 137876 703520
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106924 699712 106976 699718
rect 106924 699654 106976 699660
rect 88340 141500 88392 141506
rect 88340 141442 88392 141448
rect 84936 128308 84988 128314
rect 84936 128250 84988 128256
rect 106936 115938 106964 699654
rect 116584 656940 116636 656946
rect 116584 656882 116636 656888
rect 112444 397520 112496 397526
rect 112444 397462 112496 397468
rect 106924 115932 106976 115938
rect 106924 115874 106976 115880
rect 112456 79082 112484 397462
rect 116596 79393 116624 656882
rect 120724 616888 120776 616894
rect 120724 616830 120776 616836
rect 116676 553444 116728 553450
rect 116676 553386 116728 553392
rect 116688 79490 116716 553386
rect 118700 485104 118752 485110
rect 118700 485046 118752 485052
rect 118608 404388 118660 404394
rect 118608 404330 118660 404336
rect 118516 351960 118568 351966
rect 118516 351902 118568 351908
rect 118240 142996 118292 143002
rect 118240 142938 118292 142944
rect 118056 140140 118108 140146
rect 118056 140082 118108 140088
rect 117318 137592 117374 137601
rect 117318 137527 117374 137536
rect 117332 136746 117360 137527
rect 117320 136740 117372 136746
rect 117320 136682 117372 136688
rect 117318 136096 117374 136105
rect 117318 136031 117374 136040
rect 117332 135318 117360 136031
rect 117320 135312 117372 135318
rect 117320 135254 117372 135260
rect 117318 134600 117374 134609
rect 117318 134535 117374 134544
rect 117332 133958 117360 134535
rect 117320 133952 117372 133958
rect 117320 133894 117372 133900
rect 117412 133884 117464 133890
rect 117412 133826 117464 133832
rect 117424 133113 117452 133826
rect 117410 133104 117466 133113
rect 117410 133039 117466 133048
rect 117320 132456 117372 132462
rect 117320 132398 117372 132404
rect 117332 131617 117360 132398
rect 117318 131608 117374 131617
rect 117318 131543 117374 131552
rect 117320 131096 117372 131102
rect 117320 131038 117372 131044
rect 117332 130121 117360 131038
rect 117318 130112 117374 130121
rect 117318 130047 117374 130056
rect 117320 129736 117372 129742
rect 117320 129678 117372 129684
rect 117332 128625 117360 129678
rect 117318 128616 117374 128625
rect 117318 128551 117374 128560
rect 117320 128308 117372 128314
rect 117320 128250 117372 128256
rect 117332 127129 117360 128250
rect 117318 127120 117374 127129
rect 117318 127055 117374 127064
rect 117320 126948 117372 126954
rect 117320 126890 117372 126896
rect 117332 125633 117360 126890
rect 117318 125624 117374 125633
rect 117318 125559 117374 125568
rect 117320 124160 117372 124166
rect 117318 124128 117320 124137
rect 117372 124128 117374 124137
rect 117318 124063 117374 124072
rect 117320 122800 117372 122806
rect 117320 122742 117372 122748
rect 117332 122641 117360 122742
rect 117318 122632 117374 122641
rect 117318 122567 117374 122576
rect 117320 121440 117372 121446
rect 117320 121382 117372 121388
rect 117332 121145 117360 121382
rect 117318 121136 117374 121145
rect 117318 121071 117374 121080
rect 117320 120080 117372 120086
rect 117320 120022 117372 120028
rect 117332 119649 117360 120022
rect 117318 119640 117374 119649
rect 117318 119575 117374 119584
rect 117320 118652 117372 118658
rect 117320 118594 117372 118600
rect 117332 118153 117360 118594
rect 117318 118144 117374 118153
rect 117318 118079 117374 118088
rect 117320 117292 117372 117298
rect 117320 117234 117372 117240
rect 117332 116657 117360 117234
rect 117318 116648 117374 116657
rect 117318 116583 117374 116592
rect 117320 115932 117372 115938
rect 117320 115874 117372 115880
rect 117332 115161 117360 115874
rect 117318 115152 117374 115161
rect 117318 115087 117374 115096
rect 118068 113665 118096 140082
rect 118148 139596 118200 139602
rect 118148 139538 118200 139544
rect 118054 113656 118110 113665
rect 118054 113591 118110 113600
rect 118160 91225 118188 139538
rect 118252 92721 118280 142938
rect 118424 141568 118476 141574
rect 118424 141510 118476 141516
rect 118332 139528 118384 139534
rect 118332 139470 118384 139476
rect 118238 92712 118294 92721
rect 118238 92647 118294 92656
rect 118146 91216 118202 91225
rect 118146 91151 118202 91160
rect 118344 88233 118372 139470
rect 118436 89729 118464 141510
rect 118528 94217 118556 351902
rect 118620 95713 118648 404330
rect 118712 103193 118740 485046
rect 119344 187740 119396 187746
rect 119344 187682 119396 187688
rect 119252 147008 119304 147014
rect 119252 146950 119304 146956
rect 118976 145648 119028 145654
rect 118976 145590 119028 145596
rect 118884 141432 118936 141438
rect 118884 141374 118936 141380
rect 118792 140072 118844 140078
rect 118792 140014 118844 140020
rect 118804 104689 118832 140014
rect 118896 106185 118924 141374
rect 118988 110673 119016 145590
rect 119068 144220 119120 144226
rect 119068 144162 119120 144168
rect 118974 110664 119030 110673
rect 118974 110599 119030 110608
rect 119080 109177 119108 144162
rect 119160 142860 119212 142866
rect 119160 142802 119212 142808
rect 119066 109168 119122 109177
rect 119066 109103 119122 109112
rect 119172 107681 119200 142802
rect 119264 112169 119292 146950
rect 119250 112160 119306 112169
rect 119250 112095 119306 112104
rect 119158 107672 119214 107681
rect 119158 107607 119214 107616
rect 118882 106176 118938 106185
rect 118882 106111 118938 106120
rect 118790 104680 118846 104689
rect 118790 104615 118846 104624
rect 118698 103184 118754 103193
rect 118698 103119 118754 103128
rect 118606 95704 118662 95713
rect 118606 95639 118662 95648
rect 118514 94208 118570 94217
rect 118514 94143 118570 94152
rect 118422 89720 118478 89729
rect 118422 89655 118478 89664
rect 118330 88224 118386 88233
rect 118330 88159 118386 88168
rect 118514 86728 118570 86737
rect 118514 86663 118570 86672
rect 118422 83736 118478 83745
rect 118422 83671 118478 83680
rect 116676 79484 116728 79490
rect 116676 79426 116728 79432
rect 116582 79384 116638 79393
rect 116582 79319 116638 79328
rect 112444 79076 112496 79082
rect 112444 79018 112496 79024
rect 84844 78940 84896 78946
rect 84844 78882 84896 78888
rect 96620 78124 96672 78130
rect 96620 78066 96672 78072
rect 78680 78056 78732 78062
rect 78680 77998 78732 78004
rect 10324 77988 10376 77994
rect 10324 77930 10376 77936
rect 9036 71664 9088 71670
rect 9036 71606 9088 71612
rect 8312 16546 8800 16574
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 8772 480 8800 16546
rect 9956 3800 10008 3806
rect 9956 3742 10008 3748
rect 9968 480 9996 3742
rect 10336 3602 10364 77930
rect 67640 76764 67692 76770
rect 67640 76706 67692 76712
rect 59360 76696 59412 76702
rect 59360 76638 59412 76644
rect 34520 76628 34572 76634
rect 34520 76570 34572 76576
rect 11060 76560 11112 76566
rect 11060 76502 11112 76508
rect 11072 3602 11100 76502
rect 31760 73908 31812 73914
rect 31760 73850 31812 73856
rect 27618 72584 27674 72593
rect 27618 72519 27674 72528
rect 11150 35184 11206 35193
rect 11150 35119 11206 35128
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 11164 480 11192 35119
rect 27632 16574 27660 72519
rect 31772 16574 31800 73850
rect 27632 16546 27752 16574
rect 31772 16546 31984 16574
rect 20168 10396 20220 10402
rect 20168 10338 20220 10344
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 11992 354 12020 3538
rect 13556 480 13584 3538
rect 14752 480 14780 8910
rect 15936 7608 15988 7614
rect 15936 7550 15988 7556
rect 15948 480 15976 7550
rect 19432 4956 19484 4962
rect 19432 4898 19484 4904
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 17052 480 17080 3606
rect 18248 480 18276 4762
rect 19444 480 19472 4898
rect 12318 354 12430 480
rect 11992 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20180 354 20208 10338
rect 26514 6352 26570 6361
rect 26514 6287 26570 6296
rect 25318 6216 25374 6225
rect 24216 6180 24268 6186
rect 25318 6151 25374 6160
rect 24216 6122 24268 6128
rect 23020 5024 23072 5030
rect 23020 4966 23072 4972
rect 21824 4888 21876 4894
rect 21824 4830 21876 4836
rect 21836 480 21864 4830
rect 23032 480 23060 4966
rect 24228 480 24256 6122
rect 25332 480 25360 6151
rect 26528 480 26556 6287
rect 27724 480 27752 16546
rect 28908 7676 28960 7682
rect 28908 7618 28960 7624
rect 28920 480 28948 7618
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 30104 6248 30156 6254
rect 30104 6190 30156 6196
rect 30116 480 30144 6190
rect 31312 480 31340 6258
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 33600 6384 33652 6390
rect 33600 6326 33652 6332
rect 33612 480 33640 6326
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 76570
rect 46938 75304 46994 75313
rect 46938 75239 46994 75248
rect 41420 73976 41472 73982
rect 41420 73918 41472 73924
rect 41432 16574 41460 73918
rect 45560 36576 45612 36582
rect 45560 36518 45612 36524
rect 45572 16574 45600 36518
rect 46952 16574 46980 75239
rect 53840 75200 53892 75206
rect 53840 75142 53892 75148
rect 51080 74044 51132 74050
rect 51080 73986 51132 73992
rect 41432 16546 41920 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 35992 15904 36044 15910
rect 35992 15846 36044 15852
rect 36004 480 36032 15846
rect 40684 6588 40736 6594
rect 40684 6530 40736 6536
rect 38384 6520 38436 6526
rect 38384 6462 38436 6468
rect 37188 6452 37240 6458
rect 37188 6394 37240 6400
rect 37200 480 37228 6394
rect 38396 480 38424 6462
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 39592 480 39620 3674
rect 40696 480 40724 6530
rect 41892 480 41920 16546
rect 43076 9104 43128 9110
rect 43076 9046 43128 9052
rect 43088 480 43116 9046
rect 45466 8936 45522 8945
rect 45466 8871 45522 8880
rect 44270 7576 44326 7585
rect 44270 7511 44326 7520
rect 44284 480 44312 7511
rect 45480 480 45508 8871
rect 46676 480 46704 16546
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 50160 7744 50212 7750
rect 48962 7712 49018 7721
rect 50160 7686 50212 7692
rect 48962 7647 49018 7656
rect 48976 480 49004 7647
rect 50172 480 50200 7686
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 73986
rect 53852 16574 53880 75142
rect 57980 74112 58032 74118
rect 57980 74054 58032 74060
rect 57992 16574 58020 74054
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 53748 9036 53800 9042
rect 53748 8978 53800 8984
rect 52552 7812 52604 7818
rect 52552 7754 52604 7760
rect 52564 480 52592 7754
rect 53760 480 53788 8978
rect 54956 480 54984 16546
rect 56784 10328 56836 10334
rect 56784 10270 56836 10276
rect 56048 5092 56100 5098
rect 56048 5034 56100 5040
rect 56060 480 56088 5034
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 10270
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 76638
rect 64878 73808 64934 73817
rect 64878 73743 64934 73752
rect 60738 22672 60794 22681
rect 60738 22607 60794 22616
rect 60752 16574 60780 22607
rect 64892 16574 64920 73743
rect 60752 16546 60872 16574
rect 64892 16546 65104 16574
rect 60844 480 60872 16546
rect 64326 7984 64382 7993
rect 64326 7919 64382 7928
rect 63222 7848 63278 7857
rect 63222 7783 63278 7792
rect 62028 3868 62080 3874
rect 62028 3810 62080 3816
rect 62040 480 62068 3810
rect 63236 480 63264 7783
rect 64340 480 64368 7919
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66720 7880 66772 7886
rect 66720 7822 66772 7828
rect 66732 480 66760 7822
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 76706
rect 75920 75268 75972 75274
rect 75920 75210 75972 75216
rect 71780 72684 71832 72690
rect 71780 72626 71832 72632
rect 71792 16574 71820 72626
rect 71792 16546 72648 16574
rect 71504 10464 71556 10470
rect 71504 10406 71556 10412
rect 70308 9172 70360 9178
rect 70308 9114 70360 9120
rect 69112 3936 69164 3942
rect 69112 3878 69164 3884
rect 69124 480 69152 3878
rect 70320 480 70348 9114
rect 71516 480 71544 10406
rect 72620 480 72648 16546
rect 75000 10532 75052 10538
rect 75000 10474 75052 10480
rect 73804 9240 73856 9246
rect 73804 9182 73856 9188
rect 73816 480 73844 9182
rect 75012 480 75040 10474
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 75210
rect 78692 16574 78720 77998
rect 95882 77888 95938 77897
rect 95882 77823 95938 77832
rect 91100 76968 91152 76974
rect 91100 76910 91152 76916
rect 85580 76900 85632 76906
rect 85580 76842 85632 76848
rect 84200 76832 84252 76838
rect 84200 76774 84252 76780
rect 80058 75440 80114 75449
rect 80058 75375 80114 75384
rect 80072 16574 80100 75375
rect 82820 72548 82872 72554
rect 82820 72490 82872 72496
rect 82832 16574 82860 72490
rect 78692 16546 79272 16574
rect 80072 16546 80928 16574
rect 82832 16546 83320 16574
rect 78126 10296 78182 10305
rect 78126 10231 78182 10240
rect 77392 9308 77444 9314
rect 77392 9250 77444 9256
rect 77404 480 77432 9250
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78140 354 78168 10231
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 79244 354 79272 16546
rect 80900 480 80928 16546
rect 82084 9376 82136 9382
rect 82084 9318 82136 9324
rect 82096 480 82124 9318
rect 83292 480 83320 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 76774
rect 85592 16574 85620 76842
rect 89720 74248 89772 74254
rect 89720 74190 89772 74196
rect 86960 74180 87012 74186
rect 86960 74122 87012 74128
rect 86972 16574 87000 74122
rect 89732 16574 89760 74190
rect 91112 16574 91140 76910
rect 93860 74316 93912 74322
rect 93860 74258 93912 74264
rect 93872 16574 93900 74258
rect 85592 16546 85712 16574
rect 86972 16546 87552 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 93872 16546 94728 16574
rect 85684 480 85712 16546
rect 86868 4004 86920 4010
rect 86868 3946 86920 3952
rect 86880 480 86908 3946
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87524 354 87552 16546
rect 89168 10600 89220 10606
rect 89168 10542 89220 10548
rect 88890 6488 88946 6497
rect 88890 6423 88946 6432
rect 88904 3806 88932 6423
rect 88892 3800 88944 3806
rect 88892 3742 88944 3748
rect 89180 480 89208 10542
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 92480 10668 92532 10674
rect 92480 10610 92532 10616
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 10610
rect 93952 3800 94004 3806
rect 93952 3742 94004 3748
rect 93964 480 93992 3742
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94700 354 94728 16546
rect 95790 10432 95846 10441
rect 95896 10402 95924 77823
rect 96632 16574 96660 78066
rect 104900 77036 104952 77042
rect 104900 76978 104952 76984
rect 97998 72720 98054 72729
rect 97998 72655 98054 72664
rect 98012 16574 98040 72655
rect 102140 72616 102192 72622
rect 102140 72558 102192 72564
rect 99380 40724 99432 40730
rect 99380 40666 99432 40672
rect 99392 16574 99420 40666
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 95790 10367 95846 10376
rect 95884 10396 95936 10402
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 10367
rect 95884 10338 95936 10344
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 102152 6914 102180 72558
rect 102232 58676 102284 58682
rect 102232 58618 102284 58624
rect 102244 16574 102272 58618
rect 104912 16574 104940 76978
rect 115938 76528 115994 76537
rect 115938 76463 115994 76472
rect 114560 75404 114612 75410
rect 114560 75346 114612 75352
rect 110420 71052 110472 71058
rect 110420 70994 110472 71000
rect 102244 16546 103376 16574
rect 104912 16546 105768 16574
rect 102152 6886 102272 6914
rect 101034 3360 101090 3369
rect 101034 3295 101090 3304
rect 101048 480 101076 3295
rect 102244 480 102272 6886
rect 103348 480 103376 16546
rect 104532 5160 104584 5166
rect 104532 5102 104584 5108
rect 104544 480 104572 5102
rect 105740 480 105768 16546
rect 106464 10396 106516 10402
rect 106464 10338 106516 10344
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 10338
rect 109316 9444 109368 9450
rect 109316 9386 109368 9392
rect 108120 5228 108172 5234
rect 108120 5170 108172 5176
rect 108132 480 108160 5170
rect 109328 480 109356 9386
rect 110432 3398 110460 70994
rect 114572 16574 114600 75346
rect 115952 16574 115980 76463
rect 117320 60036 117372 60042
rect 117320 59978 117372 59984
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 114006 11656 114062 11665
rect 114006 11591 114062 11600
rect 112352 10736 112404 10742
rect 112352 10678 112404 10684
rect 110512 5296 110564 5302
rect 110512 5238 110564 5244
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 5238
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 10678
rect 114020 480 114048 11591
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 59978
rect 118436 46918 118464 83671
rect 118528 75886 118556 86663
rect 118606 85232 118662 85241
rect 118606 85167 118662 85176
rect 118620 80617 118648 85167
rect 118606 80608 118662 80617
rect 118606 80543 118662 80552
rect 119356 78441 119384 187682
rect 119436 136672 119488 136678
rect 119436 136614 119488 136620
rect 119448 79626 119476 136614
rect 120736 102105 120764 616830
rect 120816 563100 120868 563106
rect 120816 563042 120868 563048
rect 120722 102096 120778 102105
rect 120722 102031 120778 102040
rect 120828 100745 120856 563042
rect 120908 510672 120960 510678
rect 120908 510614 120960 510620
rect 120814 100736 120870 100745
rect 120814 100671 120870 100680
rect 120920 98705 120948 510614
rect 121000 456816 121052 456822
rect 121000 456758 121052 456764
rect 120906 98696 120962 98705
rect 120906 98631 120962 98640
rect 121012 97209 121040 456758
rect 121092 345092 121144 345098
rect 121092 345034 121144 345040
rect 120998 97200 121054 97209
rect 120998 97135 121054 97144
rect 120632 84244 120684 84250
rect 120632 84186 120684 84192
rect 119436 79620 119488 79626
rect 119436 79562 119488 79568
rect 120644 79558 120672 84186
rect 120722 81696 120778 81705
rect 120722 81631 120778 81640
rect 120632 79552 120684 79558
rect 120632 79494 120684 79500
rect 119342 78432 119398 78441
rect 119342 78367 119398 78376
rect 118700 78192 118752 78198
rect 118700 78134 118752 78140
rect 118516 75880 118568 75886
rect 118516 75822 118568 75828
rect 118424 46912 118476 46918
rect 118424 46854 118476 46860
rect 118712 16574 118740 78134
rect 120736 22778 120764 81631
rect 121104 79898 121132 345034
rect 146944 298172 146996 298178
rect 146944 298114 146996 298120
rect 122104 244316 122156 244322
rect 122104 244258 122156 244264
rect 122116 139602 122144 244258
rect 122196 165640 122248 165646
rect 122196 165582 122248 165588
rect 122104 139596 122156 139602
rect 122104 139538 122156 139544
rect 122208 139534 122236 165582
rect 146956 143002 146984 298114
rect 147036 205692 147088 205698
rect 147036 205634 147088 205640
rect 146944 142996 146996 143002
rect 146944 142938 146996 142944
rect 147048 141574 147076 205634
rect 147036 141568 147088 141574
rect 147036 141510 147088 141516
rect 153212 140214 153240 702406
rect 153200 140208 153252 140214
rect 153200 140150 153252 140156
rect 169772 140146 169800 702406
rect 192484 700664 192536 700670
rect 192484 700606 192536 700612
rect 190460 700324 190512 700330
rect 190460 700266 190512 700272
rect 189724 462392 189776 462398
rect 189724 462334 189776 462340
rect 189080 409896 189132 409902
rect 189080 409838 189132 409844
rect 185584 305040 185636 305046
rect 185584 304982 185636 304988
rect 185596 140554 185624 304982
rect 185584 140548 185636 140554
rect 185584 140490 185636 140496
rect 169760 140140 169812 140146
rect 169760 140082 169812 140088
rect 122196 139528 122248 139534
rect 122196 139470 122248 139476
rect 189092 121446 189120 409838
rect 189264 201544 189316 201550
rect 189264 201486 189316 201492
rect 189172 129804 189224 129810
rect 189172 129746 189224 129752
rect 189080 121440 189132 121446
rect 189080 121382 189132 121388
rect 189080 80776 189132 80782
rect 189080 80718 189132 80724
rect 188988 80708 189040 80714
rect 188988 80650 189040 80656
rect 188896 80096 188948 80102
rect 127084 80034 127296 80050
rect 127072 80028 127308 80034
rect 127124 80022 127256 80028
rect 127072 79970 127124 79976
rect 127256 79970 127308 79976
rect 130200 80028 130252 80034
rect 130200 79970 130252 79976
rect 130304 80022 130640 80050
rect 188896 80038 188948 80044
rect 127164 79960 127216 79966
rect 127164 79902 127216 79908
rect 129924 79960 129976 79966
rect 129924 79902 129976 79908
rect 130106 79928 130162 79937
rect 121092 79892 121144 79898
rect 121092 79834 121144 79840
rect 126888 79824 126940 79830
rect 126888 79766 126940 79772
rect 126336 79688 126388 79694
rect 126336 79630 126388 79636
rect 122104 78668 122156 78674
rect 122104 78610 122156 78616
rect 120724 22772 120776 22778
rect 120724 22714 120776 22720
rect 120080 19984 120132 19990
rect 120080 19926 120132 19932
rect 120092 16574 120120 19926
rect 118712 16546 118832 16574
rect 120092 16546 120672 16574
rect 118804 480 118832 16546
rect 119894 9072 119950 9081
rect 119894 9007 119950 9016
rect 119908 480 119936 9007
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122116 9110 122144 78610
rect 124862 78024 124918 78033
rect 124862 77959 124918 77968
rect 124220 62144 124272 62150
rect 124220 62086 124272 62092
rect 124232 16574 124260 62086
rect 124232 16546 124720 16574
rect 122104 9104 122156 9110
rect 122104 9046 122156 9052
rect 123484 7948 123536 7954
rect 123484 7890 123536 7896
rect 122288 5364 122340 5370
rect 122288 5306 122340 5312
rect 122300 480 122328 5306
rect 123496 480 123524 7890
rect 124692 480 124720 16546
rect 124876 15910 124904 77959
rect 126244 77308 126296 77314
rect 126244 77250 126296 77256
rect 124864 15904 124916 15910
rect 124864 15846 124916 15852
rect 125876 4072 125928 4078
rect 125876 4014 125928 4020
rect 125888 480 125916 4014
rect 126256 3534 126284 77250
rect 126348 7682 126376 79630
rect 126900 75177 126928 79766
rect 126980 77240 127032 77246
rect 126980 77182 127032 77188
rect 126886 75168 126942 75177
rect 126886 75103 126942 75112
rect 126992 11762 127020 77182
rect 127176 76566 127204 79902
rect 129464 79892 129516 79898
rect 129464 79834 129516 79840
rect 129556 79892 129608 79898
rect 129556 79834 129608 79840
rect 127624 79620 127676 79626
rect 127624 79562 127676 79568
rect 127636 79490 127664 79562
rect 129476 79558 129504 79834
rect 129372 79552 129424 79558
rect 129372 79494 129424 79500
rect 129464 79552 129516 79558
rect 129464 79494 129516 79500
rect 127624 79484 127676 79490
rect 127624 79426 127676 79432
rect 129384 79218 129412 79494
rect 129372 79212 129424 79218
rect 129372 79154 129424 79160
rect 129372 78872 129424 78878
rect 129372 78814 129424 78820
rect 127716 78260 127768 78266
rect 127716 78202 127768 78208
rect 127164 76560 127216 76566
rect 127164 76502 127216 76508
rect 127072 75472 127124 75478
rect 127072 75414 127124 75420
rect 126980 11756 127032 11762
rect 126980 11698 127032 11704
rect 126336 7676 126388 7682
rect 126336 7618 126388 7624
rect 127084 6914 127112 75414
rect 127624 73228 127676 73234
rect 127624 73170 127676 73176
rect 126992 6886 127112 6914
rect 126244 3528 126296 3534
rect 126244 3470 126296 3476
rect 126992 480 127020 6886
rect 127636 3466 127664 73170
rect 127728 62150 127756 78202
rect 129004 77852 129056 77858
rect 129004 77794 129056 77800
rect 128360 77716 128412 77722
rect 128360 77658 128412 77664
rect 127716 62144 127768 62150
rect 127716 62086 127768 62092
rect 128372 16574 128400 77658
rect 128372 16546 128952 16574
rect 128176 11756 128228 11762
rect 128176 11698 128228 11704
rect 127624 3460 127676 3466
rect 127624 3402 127676 3408
rect 128188 480 128216 11698
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 129016 3874 129044 77794
rect 129188 77784 129240 77790
rect 129188 77726 129240 77732
rect 129096 75948 129148 75954
rect 129096 75890 129148 75896
rect 129004 3868 129056 3874
rect 129004 3810 129056 3816
rect 129108 3738 129136 75890
rect 129200 5302 129228 77726
rect 129280 77444 129332 77450
rect 129280 77386 129332 77392
rect 129188 5296 129240 5302
rect 129188 5238 129240 5244
rect 129292 4962 129320 77386
rect 129384 36582 129412 78814
rect 129464 78328 129516 78334
rect 129464 78270 129516 78276
rect 129476 60042 129504 78270
rect 129568 77994 129596 79834
rect 129556 77988 129608 77994
rect 129556 77930 129608 77936
rect 129646 77752 129702 77761
rect 129646 77687 129702 77696
rect 129464 60036 129516 60042
rect 129464 59978 129516 59984
rect 129372 36576 129424 36582
rect 129372 36518 129424 36524
rect 129660 22846 129688 77687
rect 129832 77648 129884 77654
rect 129832 77590 129884 77596
rect 129844 72690 129872 77590
rect 129832 72684 129884 72690
rect 129832 72626 129884 72632
rect 129936 66910 129964 79902
rect 130106 79863 130162 79872
rect 130016 79008 130068 79014
rect 130016 78950 130068 78956
rect 130028 69698 130056 78950
rect 130016 69692 130068 69698
rect 130016 69634 130068 69640
rect 129924 66904 129976 66910
rect 129924 66846 129976 66852
rect 130120 61402 130148 79863
rect 130212 79286 130240 79970
rect 130200 79280 130252 79286
rect 130200 79222 130252 79228
rect 130304 73234 130332 80022
rect 130718 79948 130746 80036
rect 130810 79966 130838 80036
rect 130580 79920 130746 79948
rect 130798 79960 130850 79966
rect 130384 77376 130436 77382
rect 130384 77318 130436 77324
rect 130292 73228 130344 73234
rect 130292 73170 130344 73176
rect 130200 72752 130252 72758
rect 130200 72694 130252 72700
rect 130108 61396 130160 61402
rect 130108 61338 130160 61344
rect 129648 22840 129700 22846
rect 129648 22782 129700 22788
rect 130212 6914 130240 72694
rect 130396 10674 130424 77318
rect 130580 77314 130608 79920
rect 130798 79902 130850 79908
rect 130902 79744 130930 80036
rect 130994 79966 131022 80036
rect 131086 79971 131114 80036
rect 130982 79960 131034 79966
rect 130982 79902 131034 79908
rect 131072 79962 131128 79971
rect 131072 79897 131128 79906
rect 131178 79830 131206 80036
rect 131270 79898 131298 80036
rect 131258 79892 131310 79898
rect 131258 79834 131310 79840
rect 131362 79830 131390 80036
rect 131454 79971 131482 80036
rect 131440 79962 131496 79971
rect 131546 79966 131574 80036
rect 131440 79897 131496 79906
rect 131534 79960 131586 79966
rect 131534 79902 131586 79908
rect 131166 79824 131218 79830
rect 131166 79766 131218 79772
rect 131350 79824 131402 79830
rect 131638 79778 131666 80036
rect 131730 79898 131758 80036
rect 131822 79971 131850 80036
rect 131808 79962 131864 79971
rect 131718 79892 131770 79898
rect 131808 79897 131864 79906
rect 131914 79898 131942 80036
rect 132006 79966 132034 80036
rect 131994 79960 132046 79966
rect 131994 79902 132046 79908
rect 131718 79834 131770 79840
rect 131902 79892 131954 79898
rect 131902 79834 131954 79840
rect 132098 79812 132126 80036
rect 132190 79971 132218 80036
rect 132176 79962 132232 79971
rect 132176 79897 132232 79906
rect 132282 79898 132310 80036
rect 132374 79971 132402 80036
rect 132360 79962 132416 79971
rect 132270 79892 132322 79898
rect 132360 79897 132416 79906
rect 132270 79834 132322 79840
rect 131350 79766 131402 79772
rect 130856 79716 130930 79744
rect 131028 79756 131080 79762
rect 130856 79014 130884 79716
rect 131028 79698 131080 79704
rect 131592 79750 131666 79778
rect 131762 79792 131818 79801
rect 130844 79008 130896 79014
rect 130844 78950 130896 78956
rect 130844 78736 130896 78742
rect 130844 78678 130896 78684
rect 130660 78464 130712 78470
rect 130660 78406 130712 78412
rect 130568 77308 130620 77314
rect 130568 77250 130620 77256
rect 130476 72684 130528 72690
rect 130476 72626 130528 72632
rect 130488 40730 130516 72626
rect 130672 70394 130700 78406
rect 130752 77580 130804 77586
rect 130752 77522 130804 77528
rect 130764 72593 130792 77522
rect 130750 72584 130806 72593
rect 130750 72519 130806 72528
rect 130580 70366 130700 70394
rect 130580 58682 130608 70366
rect 130856 70242 130884 78678
rect 131040 77217 131068 79698
rect 131120 79688 131172 79694
rect 131592 79676 131620 79750
rect 132052 79784 132126 79812
rect 132222 79792 132278 79801
rect 131762 79727 131818 79736
rect 131856 79756 131908 79762
rect 131120 79630 131172 79636
rect 131316 79648 131620 79676
rect 131026 77208 131082 77217
rect 131026 77143 131082 77152
rect 130936 75540 130988 75546
rect 130936 75482 130988 75488
rect 130948 72962 130976 75482
rect 131132 73273 131160 79630
rect 131316 76616 131344 79648
rect 131394 78160 131450 78169
rect 131394 78095 131450 78104
rect 131224 76588 131344 76616
rect 131118 73264 131174 73273
rect 131118 73199 131174 73208
rect 130936 72956 130988 72962
rect 130936 72898 130988 72904
rect 130844 70236 130896 70242
rect 130844 70178 130896 70184
rect 130568 58676 130620 58682
rect 130568 58618 130620 58624
rect 130476 40724 130528 40730
rect 130476 40666 130528 40672
rect 130384 10668 130436 10674
rect 130384 10610 130436 10616
rect 130212 6886 130608 6914
rect 129280 4956 129332 4962
rect 129280 4898 129332 4904
rect 129096 3732 129148 3738
rect 129096 3674 129148 3680
rect 130580 480 130608 6886
rect 131224 3602 131252 76588
rect 131304 75608 131356 75614
rect 131304 75550 131356 75556
rect 131316 75274 131344 75550
rect 131304 75268 131356 75274
rect 131304 75210 131356 75216
rect 131304 75132 131356 75138
rect 131304 75074 131356 75080
rect 131316 4894 131344 75074
rect 131408 5030 131436 78095
rect 131776 78010 131804 79727
rect 131856 79698 131908 79704
rect 131488 77988 131540 77994
rect 131488 77930 131540 77936
rect 131592 77982 131804 78010
rect 131500 76514 131528 77930
rect 131592 77160 131620 77982
rect 131672 77920 131724 77926
rect 131672 77862 131724 77868
rect 131684 77228 131712 77862
rect 131868 77602 131896 79698
rect 131948 79688 132000 79694
rect 131948 79630 132000 79636
rect 131960 77926 131988 79630
rect 131948 77920 132000 77926
rect 131948 77862 132000 77868
rect 131868 77574 131988 77602
rect 131856 77512 131908 77518
rect 131856 77454 131908 77460
rect 131684 77200 131804 77228
rect 131592 77132 131712 77160
rect 131500 76486 131620 76514
rect 131488 76424 131540 76430
rect 131488 76366 131540 76372
rect 131396 5024 131448 5030
rect 131396 4966 131448 4972
rect 131304 4888 131356 4894
rect 131304 4830 131356 4836
rect 131500 4826 131528 76366
rect 131592 6186 131620 76486
rect 131684 7614 131712 77132
rect 131776 8974 131804 77200
rect 131868 76770 131896 77454
rect 131856 76764 131908 76770
rect 131856 76706 131908 76712
rect 131764 8968 131816 8974
rect 131764 8910 131816 8916
rect 131672 7608 131724 7614
rect 131672 7550 131724 7556
rect 131580 6180 131632 6186
rect 131580 6122 131632 6128
rect 131488 4820 131540 4826
rect 131488 4762 131540 4768
rect 131960 3670 131988 77574
rect 132052 77450 132080 79784
rect 132144 79736 132222 79744
rect 132466 79744 132494 80036
rect 132558 79830 132586 80036
rect 132546 79824 132598 79830
rect 132650 79812 132678 80036
rect 132742 79937 132770 80036
rect 132728 79928 132784 79937
rect 132834 79898 132862 80036
rect 132926 79971 132954 80036
rect 132912 79962 132968 79971
rect 132728 79863 132784 79872
rect 132822 79892 132874 79898
rect 132912 79897 132968 79906
rect 132822 79834 132874 79840
rect 132650 79801 132724 79812
rect 132650 79792 132738 79801
rect 132650 79784 132682 79792
rect 132546 79766 132598 79772
rect 132144 79727 132278 79736
rect 132144 79716 132264 79727
rect 132420 79716 132494 79744
rect 132682 79727 132738 79736
rect 132144 77586 132172 79716
rect 132224 79620 132276 79626
rect 132224 79562 132276 79568
rect 132132 77580 132184 77586
rect 132132 77522 132184 77528
rect 132040 77444 132092 77450
rect 132040 77386 132092 77392
rect 132132 77444 132184 77450
rect 132132 77386 132184 77392
rect 132144 73914 132172 77386
rect 132236 76430 132264 79562
rect 132420 77994 132448 79716
rect 132592 79688 132644 79694
rect 132592 79630 132644 79636
rect 132684 79688 132736 79694
rect 132684 79630 132736 79636
rect 132868 79688 132920 79694
rect 133018 79676 133046 80036
rect 133110 79744 133138 80036
rect 133202 79898 133230 80036
rect 133294 79971 133322 80036
rect 133280 79962 133336 79971
rect 133386 79966 133414 80036
rect 133190 79892 133242 79898
rect 133280 79897 133336 79906
rect 133374 79960 133426 79966
rect 133478 79937 133506 80036
rect 133570 79966 133598 80036
rect 133662 79971 133690 80036
rect 133558 79960 133610 79966
rect 133374 79902 133426 79908
rect 133464 79928 133520 79937
rect 133558 79902 133610 79908
rect 133648 79962 133704 79971
rect 133754 79966 133782 80036
rect 133846 79966 133874 80036
rect 133648 79897 133704 79906
rect 133742 79960 133794 79966
rect 133742 79902 133794 79908
rect 133834 79960 133886 79966
rect 133834 79902 133886 79908
rect 133464 79863 133520 79872
rect 133190 79834 133242 79840
rect 133696 79824 133748 79830
rect 133234 79792 133290 79801
rect 133110 79716 133184 79744
rect 133234 79727 133290 79736
rect 133418 79792 133474 79801
rect 133602 79792 133658 79801
rect 133418 79727 133474 79736
rect 133512 79756 133564 79762
rect 133018 79648 133092 79676
rect 132868 79630 132920 79636
rect 132500 79620 132552 79626
rect 132500 79562 132552 79568
rect 132408 77988 132460 77994
rect 132408 77930 132460 77936
rect 132408 77308 132460 77314
rect 132408 77250 132460 77256
rect 132224 76424 132276 76430
rect 132224 76366 132276 76372
rect 132420 75313 132448 77250
rect 132406 75304 132462 75313
rect 132406 75239 132462 75248
rect 132512 75138 132540 79562
rect 132604 75857 132632 79630
rect 132696 79286 132724 79630
rect 132684 79280 132736 79286
rect 132684 79222 132736 79228
rect 132880 78248 132908 79630
rect 132880 78220 133000 78248
rect 132866 78160 132922 78169
rect 132866 78095 132922 78104
rect 132684 76560 132736 76566
rect 132684 76502 132736 76508
rect 132590 75848 132646 75857
rect 132590 75783 132646 75792
rect 132500 75132 132552 75138
rect 132500 75074 132552 75080
rect 132132 73908 132184 73914
rect 132132 73850 132184 73856
rect 132696 6594 132724 76502
rect 132776 73704 132828 73710
rect 132776 73646 132828 73652
rect 132684 6588 132736 6594
rect 132684 6530 132736 6536
rect 132788 6458 132816 73646
rect 132776 6452 132828 6458
rect 132776 6394 132828 6400
rect 132880 6254 132908 78095
rect 132972 6390 133000 78220
rect 133064 76752 133092 79648
rect 133156 77450 133184 79716
rect 133144 77444 133196 77450
rect 133144 77386 133196 77392
rect 133064 76724 133184 76752
rect 133052 76628 133104 76634
rect 133052 76570 133104 76576
rect 133064 6526 133092 76570
rect 133052 6520 133104 6526
rect 133052 6462 133104 6468
rect 132960 6384 133012 6390
rect 132960 6326 133012 6332
rect 133156 6322 133184 76724
rect 133248 76498 133276 79727
rect 133328 79688 133380 79694
rect 133328 79630 133380 79636
rect 133340 78033 133368 79630
rect 133326 78024 133382 78033
rect 133326 77959 133382 77968
rect 133236 76492 133288 76498
rect 133236 76434 133288 76440
rect 133432 73710 133460 79727
rect 133938 79778 133966 80036
rect 134030 79971 134058 80036
rect 134016 79962 134072 79971
rect 134016 79897 134072 79906
rect 134122 79812 134150 80036
rect 134214 79966 134242 80036
rect 134202 79960 134254 79966
rect 134202 79902 134254 79908
rect 134076 79801 134150 79812
rect 133696 79766 133748 79772
rect 133602 79727 133658 79736
rect 133512 79698 133564 79704
rect 133524 76634 133552 79698
rect 133512 76628 133564 76634
rect 133512 76570 133564 76576
rect 133616 75954 133644 79727
rect 133708 76566 133736 79766
rect 133892 79750 133966 79778
rect 134062 79792 134150 79801
rect 133788 79688 133840 79694
rect 133788 79630 133840 79636
rect 133696 76560 133748 76566
rect 133696 76502 133748 76508
rect 133604 75948 133656 75954
rect 133604 75890 133656 75896
rect 133800 73982 133828 79630
rect 133892 78810 133920 79750
rect 134118 79784 134150 79792
rect 134062 79727 134118 79736
rect 134064 79688 134116 79694
rect 134064 79630 134116 79636
rect 133880 78804 133932 78810
rect 133880 78746 133932 78752
rect 133970 78704 134026 78713
rect 133970 78639 134026 78648
rect 133788 73976 133840 73982
rect 133788 73918 133840 73924
rect 133420 73704 133472 73710
rect 133420 73646 133472 73652
rect 133144 6316 133196 6322
rect 133144 6258 133196 6264
rect 132868 6248 132920 6254
rect 132868 6190 132920 6196
rect 131948 3664 132000 3670
rect 131948 3606 132000 3612
rect 131212 3596 131264 3602
rect 131212 3538 131264 3544
rect 131764 3528 131816 3534
rect 131764 3470 131816 3476
rect 131776 480 131804 3470
rect 132960 3460 133012 3466
rect 132960 3402 133012 3408
rect 132972 480 133000 3402
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133984 354 134012 78639
rect 134076 7818 134104 79630
rect 134156 79620 134208 79626
rect 134156 79562 134208 79568
rect 134168 78878 134196 79562
rect 134306 79540 134334 80036
rect 134398 79801 134426 80036
rect 134384 79792 134440 79801
rect 134384 79727 134440 79736
rect 134490 79608 134518 80036
rect 134582 79778 134610 80036
rect 134674 79898 134702 80036
rect 134662 79892 134714 79898
rect 134662 79834 134714 79840
rect 134766 79778 134794 80036
rect 134582 79750 134656 79778
rect 134260 79512 134334 79540
rect 134444 79580 134518 79608
rect 134156 78872 134208 78878
rect 134156 78814 134208 78820
rect 134260 77314 134288 79512
rect 134444 78656 134472 79580
rect 134524 79280 134576 79286
rect 134524 79222 134576 79228
rect 134352 78628 134472 78656
rect 134248 77308 134300 77314
rect 134248 77250 134300 77256
rect 134352 77160 134380 78628
rect 134432 78532 134484 78538
rect 134432 78474 134484 78480
rect 134168 77132 134380 77160
rect 134064 7812 134116 7818
rect 134064 7754 134116 7760
rect 134168 7750 134196 77132
rect 134248 75268 134300 75274
rect 134248 75210 134300 75216
rect 134260 9042 134288 75210
rect 134340 75200 134392 75206
rect 134340 75142 134392 75148
rect 134352 10334 134380 75142
rect 134340 10328 134392 10334
rect 134340 10270 134392 10276
rect 134248 9036 134300 9042
rect 134248 8978 134300 8984
rect 134156 7744 134208 7750
rect 134156 7686 134208 7692
rect 134444 5098 134472 78474
rect 134536 78266 134564 79222
rect 134524 78260 134576 78266
rect 134524 78202 134576 78208
rect 134524 77308 134576 77314
rect 134524 77250 134576 77256
rect 134536 10538 134564 77250
rect 134628 74050 134656 79750
rect 134720 79750 134794 79778
rect 134858 79778 134886 80036
rect 134950 79898 134978 80036
rect 135042 79937 135070 80036
rect 135028 79928 135084 79937
rect 134938 79892 134990 79898
rect 135134 79898 135162 80036
rect 135226 79966 135254 80036
rect 135214 79960 135266 79966
rect 135214 79902 135266 79908
rect 135028 79863 135084 79872
rect 135122 79892 135174 79898
rect 134938 79834 134990 79840
rect 135122 79834 135174 79840
rect 135318 79812 135346 80036
rect 135272 79801 135346 79812
rect 135258 79792 135346 79801
rect 134858 79750 134932 79778
rect 134720 75274 134748 79750
rect 134800 79688 134852 79694
rect 134800 79630 134852 79636
rect 134812 78538 134840 79630
rect 134800 78532 134852 78538
rect 134800 78474 134852 78480
rect 134708 75268 134760 75274
rect 134708 75210 134760 75216
rect 134904 75070 134932 79750
rect 135314 79784 135346 79792
rect 135410 79744 135438 80036
rect 135502 79937 135530 80036
rect 135488 79928 135544 79937
rect 135488 79863 135544 79872
rect 135594 79778 135622 80036
rect 135686 79801 135714 80036
rect 135258 79727 135314 79736
rect 135364 79716 135438 79744
rect 135548 79750 135622 79778
rect 135672 79792 135728 79801
rect 135076 79688 135128 79694
rect 135076 79630 135128 79636
rect 135168 79688 135220 79694
rect 135168 79630 135220 79636
rect 135088 78826 135116 79630
rect 134996 78798 135116 78826
rect 134892 75064 134944 75070
rect 134892 75006 134944 75012
rect 134996 74118 135024 78798
rect 135074 78704 135130 78713
rect 135074 78639 135130 78648
rect 135088 75206 135116 78639
rect 135180 76702 135208 79630
rect 135364 79608 135392 79716
rect 135272 79580 135392 79608
rect 135272 77858 135300 79580
rect 135444 79552 135496 79558
rect 135444 79494 135496 79500
rect 135352 79484 135404 79490
rect 135352 79426 135404 79432
rect 135364 78878 135392 79426
rect 135352 78872 135404 78878
rect 135352 78814 135404 78820
rect 135260 77852 135312 77858
rect 135260 77794 135312 77800
rect 135260 77580 135312 77586
rect 135260 77522 135312 77528
rect 135168 76696 135220 76702
rect 135168 76638 135220 76644
rect 135076 75200 135128 75206
rect 135076 75142 135128 75148
rect 134984 74112 135036 74118
rect 134984 74054 135036 74060
rect 134616 74044 134668 74050
rect 134616 73986 134668 73992
rect 135272 11762 135300 77522
rect 135456 77294 135484 79494
rect 135548 77353 135576 79750
rect 135672 79727 135728 79736
rect 135628 79688 135680 79694
rect 135628 79630 135680 79636
rect 135640 77518 135668 79630
rect 135778 79506 135806 80036
rect 135870 79898 135898 80036
rect 135962 79898 135990 80036
rect 135858 79892 135910 79898
rect 135858 79834 135910 79840
rect 135950 79892 136002 79898
rect 135950 79834 136002 79840
rect 136054 79744 136082 80036
rect 136008 79716 136082 79744
rect 135904 79620 135956 79626
rect 135904 79562 135956 79568
rect 135732 79478 135806 79506
rect 135628 77512 135680 77518
rect 135628 77454 135680 77460
rect 135364 77266 135484 77294
rect 135534 77344 135590 77353
rect 135534 77279 135590 77288
rect 135260 11756 135312 11762
rect 135260 11698 135312 11704
rect 134524 10532 134576 10538
rect 134524 10474 134576 10480
rect 135260 8152 135312 8158
rect 135260 8094 135312 8100
rect 134432 5092 134484 5098
rect 134432 5034 134484 5040
rect 135272 480 135300 8094
rect 135364 3942 135392 77266
rect 135732 77058 135760 79478
rect 135916 79121 135944 79562
rect 135902 79112 135958 79121
rect 135902 79047 135958 79056
rect 136008 78962 136036 79716
rect 136146 79676 136174 80036
rect 135548 77030 135760 77058
rect 135824 78934 136036 78962
rect 136100 79648 136174 79676
rect 135444 71800 135496 71806
rect 135444 71742 135496 71748
rect 135456 8158 135484 71742
rect 135444 8152 135496 8158
rect 135444 8094 135496 8100
rect 135548 7886 135576 77030
rect 135628 75268 135680 75274
rect 135628 75210 135680 75216
rect 135640 9246 135668 75210
rect 135720 75200 135772 75206
rect 135720 75142 135772 75148
rect 135732 9314 135760 75142
rect 135720 9308 135772 9314
rect 135720 9250 135772 9256
rect 135628 9240 135680 9246
rect 135628 9182 135680 9188
rect 135824 9178 135852 78934
rect 135996 78804 136048 78810
rect 135996 78746 136048 78752
rect 136008 73030 136036 78746
rect 135996 73024 136048 73030
rect 135996 72966 136048 72972
rect 136100 70394 136128 79648
rect 136238 79608 136266 80036
rect 136330 79676 136358 80036
rect 136422 79744 136450 80036
rect 136514 79937 136542 80036
rect 136500 79928 136556 79937
rect 136606 79898 136634 80036
rect 136698 79966 136726 80036
rect 136790 79966 136818 80036
rect 136882 79966 136910 80036
rect 136686 79960 136738 79966
rect 136686 79902 136738 79908
rect 136778 79960 136830 79966
rect 136778 79902 136830 79908
rect 136870 79960 136922 79966
rect 136870 79902 136922 79908
rect 136500 79863 136556 79872
rect 136594 79892 136646 79898
rect 136594 79834 136646 79840
rect 136824 79824 136876 79830
rect 136638 79792 136694 79801
rect 136422 79716 136496 79744
rect 136824 79766 136876 79772
rect 136638 79727 136694 79736
rect 136732 79756 136784 79762
rect 136330 79648 136404 79676
rect 136192 79580 136266 79608
rect 136192 78810 136220 79580
rect 136272 79484 136324 79490
rect 136272 79426 136324 79432
rect 136284 78849 136312 79426
rect 136270 78840 136326 78849
rect 136180 78804 136232 78810
rect 136270 78775 136326 78784
rect 136180 78746 136232 78752
rect 136178 78704 136234 78713
rect 136376 78656 136404 79648
rect 136178 78639 136234 78648
rect 136192 75614 136220 78639
rect 136284 78628 136404 78656
rect 136180 75608 136232 75614
rect 136180 75550 136232 75556
rect 136284 75274 136312 78628
rect 136364 78532 136416 78538
rect 136364 78474 136416 78480
rect 136376 76906 136404 78474
rect 136468 77314 136496 79716
rect 136548 79688 136600 79694
rect 136548 79630 136600 79636
rect 136456 77308 136508 77314
rect 136456 77250 136508 77256
rect 136364 76900 136416 76906
rect 136364 76842 136416 76848
rect 136272 75268 136324 75274
rect 136272 75210 136324 75216
rect 136560 75206 136588 79630
rect 136652 76838 136680 79727
rect 136732 79698 136784 79704
rect 136744 78713 136772 79698
rect 136730 78704 136786 78713
rect 136730 78639 136786 78648
rect 136836 78062 136864 79766
rect 136974 79676 137002 80036
rect 137066 79937 137094 80036
rect 137052 79928 137108 79937
rect 137052 79863 137108 79872
rect 137158 79801 137186 80036
rect 137144 79792 137200 79801
rect 137144 79727 137200 79736
rect 136928 79648 137002 79676
rect 137100 79688 137152 79694
rect 136824 78056 136876 78062
rect 136824 77998 136876 78004
rect 136730 77888 136786 77897
rect 136730 77823 136786 77832
rect 136744 77654 136772 77823
rect 136732 77648 136784 77654
rect 136732 77590 136784 77596
rect 136640 76832 136692 76838
rect 136640 76774 136692 76780
rect 136548 75200 136600 75206
rect 136548 75142 136600 75148
rect 136824 73228 136876 73234
rect 136824 73170 136876 73176
rect 135916 70366 136128 70394
rect 135916 10470 135944 70366
rect 136456 11756 136508 11762
rect 136456 11698 136508 11704
rect 135904 10464 135956 10470
rect 135904 10406 135956 10412
rect 135812 9172 135864 9178
rect 135812 9114 135864 9120
rect 135536 7880 135588 7886
rect 135536 7822 135588 7828
rect 135352 3936 135404 3942
rect 135352 3878 135404 3884
rect 136468 480 136496 11698
rect 136836 6914 136864 73170
rect 136928 9382 136956 79648
rect 137250 79676 137278 80036
rect 137342 79744 137370 80036
rect 137434 79812 137462 80036
rect 137526 79966 137554 80036
rect 137514 79960 137566 79966
rect 137514 79902 137566 79908
rect 137618 79812 137646 80036
rect 137434 79784 137508 79812
rect 137342 79716 137416 79744
rect 137100 79630 137152 79636
rect 137204 79648 137278 79676
rect 137008 79552 137060 79558
rect 137008 79494 137060 79500
rect 137020 10606 137048 79494
rect 137008 10600 137060 10606
rect 137008 10542 137060 10548
rect 136916 9376 136968 9382
rect 136916 9318 136968 9324
rect 136836 6886 137048 6914
rect 137020 490 137048 6886
rect 137112 3806 137140 79630
rect 137204 78538 137232 79648
rect 137284 79144 137336 79150
rect 137284 79086 137336 79092
rect 137192 78532 137244 78538
rect 137192 78474 137244 78480
rect 137296 75342 137324 79086
rect 137284 75336 137336 75342
rect 137284 75278 137336 75284
rect 137388 70394 137416 79716
rect 137480 74186 137508 79784
rect 137572 79784 137646 79812
rect 137572 74254 137600 79784
rect 137710 79744 137738 80036
rect 137802 79778 137830 80036
rect 137894 79898 137922 80036
rect 137882 79892 137934 79898
rect 137882 79834 137934 79840
rect 137986 79778 138014 80036
rect 137802 79750 137876 79778
rect 137664 79716 137738 79744
rect 137664 76974 137692 79716
rect 137744 79484 137796 79490
rect 137744 79426 137796 79432
rect 137756 78849 137784 79426
rect 137742 78840 137798 78849
rect 137742 78775 137798 78784
rect 137742 78704 137798 78713
rect 137742 78639 137798 78648
rect 137652 76968 137704 76974
rect 137652 76910 137704 76916
rect 137560 74248 137612 74254
rect 137560 74190 137612 74196
rect 137468 74180 137520 74186
rect 137468 74122 137520 74128
rect 137756 72554 137784 78639
rect 137848 77382 137876 79750
rect 137940 79750 138014 79778
rect 138078 79778 138106 80036
rect 138170 79966 138198 80036
rect 138158 79960 138210 79966
rect 138158 79902 138210 79908
rect 138262 79812 138290 80036
rect 138354 79971 138382 80036
rect 138340 79962 138396 79971
rect 138340 79897 138396 79906
rect 138262 79801 138336 79812
rect 138262 79792 138350 79801
rect 138262 79784 138294 79792
rect 138078 79750 138152 79778
rect 137836 77376 137888 77382
rect 137836 77318 137888 77324
rect 137940 74322 137968 79750
rect 138020 79688 138072 79694
rect 138020 79630 138072 79636
rect 138032 78130 138060 79630
rect 138124 78713 138152 79750
rect 138446 79778 138474 80036
rect 138538 79937 138566 80036
rect 138524 79928 138580 79937
rect 138524 79863 138580 79872
rect 138630 79812 138658 80036
rect 138294 79727 138350 79736
rect 138400 79750 138474 79778
rect 138584 79784 138658 79812
rect 138296 79688 138348 79694
rect 138296 79630 138348 79636
rect 138202 78976 138258 78985
rect 138202 78911 138258 78920
rect 138110 78704 138166 78713
rect 138110 78639 138166 78648
rect 138020 78124 138072 78130
rect 138020 78066 138072 78072
rect 138020 75948 138072 75954
rect 138020 75890 138072 75896
rect 137928 74316 137980 74322
rect 137928 74258 137980 74264
rect 137744 72548 137796 72554
rect 137744 72490 137796 72496
rect 137296 70366 137416 70394
rect 137296 4010 137324 70366
rect 138032 16574 138060 75890
rect 138032 16546 138152 16574
rect 137284 4004 137336 4010
rect 137284 3946 137336 3952
rect 137100 3800 137152 3806
rect 137100 3742 137152 3748
rect 138124 3482 138152 16546
rect 138216 5234 138244 78911
rect 138308 9450 138336 79630
rect 138400 78849 138428 79750
rect 138480 79688 138532 79694
rect 138480 79630 138532 79636
rect 138386 78840 138442 78849
rect 138386 78775 138442 78784
rect 138388 75268 138440 75274
rect 138388 75210 138440 75216
rect 138400 10742 138428 75210
rect 138388 10736 138440 10742
rect 138388 10678 138440 10684
rect 138492 10402 138520 79630
rect 138584 78962 138612 79784
rect 138722 79676 138750 80036
rect 138814 79744 138842 80036
rect 138906 79898 138934 80036
rect 138998 79937 139026 80036
rect 138984 79928 139040 79937
rect 138894 79892 138946 79898
rect 139090 79898 139118 80036
rect 138984 79863 139040 79872
rect 139078 79892 139130 79898
rect 138894 79834 138946 79840
rect 139078 79834 139130 79840
rect 138938 79792 138994 79801
rect 138814 79716 138888 79744
rect 139182 79778 139210 80036
rect 139274 79898 139302 80036
rect 139262 79892 139314 79898
rect 139262 79834 139314 79840
rect 138938 79727 138994 79736
rect 139044 79750 139210 79778
rect 138722 79648 138796 79676
rect 138584 78934 138704 78962
rect 138572 78736 138624 78742
rect 138572 78678 138624 78684
rect 138584 71058 138612 78678
rect 138676 78470 138704 78934
rect 138664 78464 138716 78470
rect 138664 78406 138716 78412
rect 138572 71052 138624 71058
rect 138572 70994 138624 71000
rect 138768 70394 138796 79648
rect 138860 77042 138888 79716
rect 138848 77036 138900 77042
rect 138848 76978 138900 76984
rect 138952 72622 138980 79727
rect 139044 77790 139072 79750
rect 139366 79744 139394 80036
rect 139320 79716 139394 79744
rect 139124 79688 139176 79694
rect 139124 79630 139176 79636
rect 139032 77784 139084 77790
rect 139032 77726 139084 77732
rect 139136 75410 139164 79630
rect 139216 79620 139268 79626
rect 139216 79562 139268 79568
rect 139228 78742 139256 79562
rect 139216 78736 139268 78742
rect 139216 78678 139268 78684
rect 139124 75404 139176 75410
rect 139124 75346 139176 75352
rect 139320 75274 139348 79716
rect 139458 79676 139486 80036
rect 139550 79966 139578 80036
rect 139642 79971 139670 80036
rect 139538 79960 139590 79966
rect 139538 79902 139590 79908
rect 139628 79962 139684 79971
rect 139628 79897 139684 79906
rect 139734 79898 139762 80036
rect 139722 79892 139774 79898
rect 139722 79834 139774 79840
rect 139826 79830 139854 80036
rect 139918 79937 139946 80036
rect 139904 79928 139960 79937
rect 139904 79863 139960 79872
rect 139814 79824 139866 79830
rect 139814 79766 139866 79772
rect 140010 79744 140038 80036
rect 140102 79898 140130 80036
rect 140194 79898 140222 80036
rect 140286 79971 140314 80036
rect 140272 79962 140328 79971
rect 140378 79966 140406 80036
rect 140470 79966 140498 80036
rect 140562 79966 140590 80036
rect 140090 79892 140142 79898
rect 140090 79834 140142 79840
rect 140182 79892 140234 79898
rect 140272 79897 140328 79906
rect 140366 79960 140418 79966
rect 140366 79902 140418 79908
rect 140458 79960 140510 79966
rect 140458 79902 140510 79908
rect 140550 79960 140602 79966
rect 140550 79902 140602 79908
rect 140654 79898 140682 80036
rect 140746 79937 140774 80036
rect 140732 79928 140788 79937
rect 140182 79834 140234 79840
rect 140642 79892 140694 79898
rect 140732 79863 140788 79872
rect 140642 79834 140694 79840
rect 140320 79824 140372 79830
rect 139964 79716 140038 79744
rect 140134 79792 140190 79801
rect 140838 79812 140866 80036
rect 140320 79766 140372 79772
rect 140594 79792 140650 79801
rect 140134 79727 140190 79736
rect 139584 79688 139636 79694
rect 139458 79648 139532 79676
rect 139400 79552 139452 79558
rect 139400 79494 139452 79500
rect 139412 78198 139440 79494
rect 139504 78713 139532 79648
rect 139584 79630 139636 79636
rect 139490 78704 139546 78713
rect 139490 78639 139546 78648
rect 139596 78334 139624 79630
rect 139964 79608 139992 79716
rect 139688 79580 139992 79608
rect 140044 79620 140096 79626
rect 139584 78328 139636 78334
rect 139584 78270 139636 78276
rect 139400 78192 139452 78198
rect 139400 78134 139452 78140
rect 139308 75268 139360 75274
rect 139308 75210 139360 75216
rect 139584 75268 139636 75274
rect 139584 75210 139636 75216
rect 138940 72616 138992 72622
rect 138940 72558 138992 72564
rect 138768 70366 138980 70394
rect 138480 10396 138532 10402
rect 138480 10338 138532 10344
rect 138296 9444 138348 9450
rect 138296 9386 138348 9392
rect 138204 5228 138256 5234
rect 138204 5170 138256 5176
rect 138952 5166 138980 70366
rect 139596 7954 139624 75210
rect 139688 19990 139716 79580
rect 140044 79562 140096 79568
rect 139768 79484 139820 79490
rect 139768 79426 139820 79432
rect 139676 19984 139728 19990
rect 139676 19926 139728 19932
rect 139584 7948 139636 7954
rect 139584 7890 139636 7896
rect 138940 5160 138992 5166
rect 138940 5102 138992 5108
rect 139780 4078 139808 79426
rect 140056 79370 140084 79562
rect 139964 79342 140084 79370
rect 139964 5370 139992 79342
rect 140148 79286 140176 79727
rect 140228 79688 140280 79694
rect 140228 79630 140280 79636
rect 140136 79280 140188 79286
rect 140136 79222 140188 79228
rect 140044 79212 140096 79218
rect 140044 79154 140096 79160
rect 140056 78946 140084 79154
rect 140136 79144 140188 79150
rect 140136 79086 140188 79092
rect 140044 78940 140096 78946
rect 140044 78882 140096 78888
rect 140044 78736 140096 78742
rect 140044 78678 140096 78684
rect 139952 5364 140004 5370
rect 139952 5306 140004 5312
rect 139768 4072 139820 4078
rect 139768 4014 139820 4020
rect 140056 3534 140084 78678
rect 140148 78470 140176 79086
rect 140136 78464 140188 78470
rect 140136 78406 140188 78412
rect 140136 78328 140188 78334
rect 140136 78270 140188 78276
rect 140044 3528 140096 3534
rect 138124 3454 138888 3482
rect 140044 3470 140096 3476
rect 140148 3466 140176 78270
rect 140240 75274 140268 79630
rect 140332 75478 140360 79766
rect 140412 79756 140464 79762
rect 140594 79727 140650 79736
rect 140792 79784 140866 79812
rect 140412 79698 140464 79704
rect 140424 77246 140452 79698
rect 140504 79552 140556 79558
rect 140504 79494 140556 79500
rect 140516 78742 140544 79494
rect 140504 78736 140556 78742
rect 140504 78678 140556 78684
rect 140412 77240 140464 77246
rect 140412 77182 140464 77188
rect 140608 75546 140636 79727
rect 140792 79626 140820 79784
rect 140930 79744 140958 80036
rect 141022 79898 141050 80036
rect 141010 79892 141062 79898
rect 141010 79834 141062 79840
rect 141114 79778 141142 80036
rect 141206 79835 141234 80036
rect 140884 79716 140958 79744
rect 141068 79750 141142 79778
rect 141192 79826 141248 79835
rect 141298 79812 141326 80036
rect 141390 79966 141418 80036
rect 141482 79966 141510 80036
rect 141378 79960 141430 79966
rect 141378 79902 141430 79908
rect 141470 79960 141522 79966
rect 141470 79902 141522 79908
rect 141298 79784 141372 79812
rect 141192 79761 141248 79770
rect 140780 79620 140832 79626
rect 140780 79562 140832 79568
rect 140780 79484 140832 79490
rect 140780 79426 140832 79432
rect 140792 77722 140820 79426
rect 140884 78334 140912 79716
rect 141068 79642 141096 79750
rect 140976 79614 141096 79642
rect 141240 79688 141292 79694
rect 141240 79630 141292 79636
rect 141148 79620 141200 79626
rect 140976 79354 141004 79614
rect 141148 79562 141200 79568
rect 141056 79552 141108 79558
rect 141056 79494 141108 79500
rect 140964 79348 141016 79354
rect 140964 79290 141016 79296
rect 140964 79212 141016 79218
rect 140964 79154 141016 79160
rect 140872 78328 140924 78334
rect 140872 78270 140924 78276
rect 140780 77716 140832 77722
rect 140780 77658 140832 77664
rect 140870 77616 140926 77625
rect 140870 77551 140872 77560
rect 140924 77551 140926 77560
rect 140872 77522 140924 77528
rect 140688 77444 140740 77450
rect 140688 77386 140740 77392
rect 140596 75540 140648 75546
rect 140596 75482 140648 75488
rect 140320 75472 140372 75478
rect 140320 75414 140372 75420
rect 140228 75268 140280 75274
rect 140228 75210 140280 75216
rect 140700 3738 140728 77386
rect 140976 4146 141004 79154
rect 140964 4140 141016 4146
rect 140964 4082 141016 4088
rect 140688 3732 140740 3738
rect 140688 3674 140740 3680
rect 141068 3602 141096 79494
rect 141056 3596 141108 3602
rect 141056 3538 141108 3544
rect 134126 354 134238 480
rect 133984 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137020 462 137232 490
rect 138860 480 138888 3454
rect 140136 3460 140188 3466
rect 140136 3402 140188 3408
rect 141160 3058 141188 79562
rect 141252 78792 141280 79630
rect 141344 79608 141372 79784
rect 141574 79744 141602 80036
rect 141666 79937 141694 80036
rect 141758 79966 141786 80036
rect 141850 79966 141878 80036
rect 141942 79966 141970 80036
rect 142034 79966 142062 80036
rect 142126 79966 142154 80036
rect 141746 79960 141798 79966
rect 141652 79928 141708 79937
rect 141746 79902 141798 79908
rect 141838 79960 141890 79966
rect 141838 79902 141890 79908
rect 141930 79960 141982 79966
rect 141930 79902 141982 79908
rect 142022 79960 142074 79966
rect 142022 79902 142074 79908
rect 142114 79960 142166 79966
rect 142114 79902 142166 79908
rect 141652 79863 141708 79872
rect 141700 79824 141752 79830
rect 142218 79778 142246 80036
rect 142310 79966 142338 80036
rect 142298 79960 142350 79966
rect 142298 79902 142350 79908
rect 142402 79898 142430 80036
rect 142494 79898 142522 80036
rect 142586 79898 142614 80036
rect 142678 79937 142706 80036
rect 142770 79966 142798 80036
rect 142758 79960 142810 79966
rect 142664 79928 142720 79937
rect 142390 79892 142442 79898
rect 142390 79834 142442 79840
rect 142482 79892 142534 79898
rect 142482 79834 142534 79840
rect 142574 79892 142626 79898
rect 142758 79902 142810 79908
rect 142664 79863 142720 79872
rect 142574 79834 142626 79840
rect 142862 79812 142890 80036
rect 142954 79966 142982 80036
rect 143046 79966 143074 80036
rect 142942 79960 142994 79966
rect 142942 79902 142994 79908
rect 143034 79960 143086 79966
rect 143034 79902 143086 79908
rect 142988 79824 143040 79830
rect 142862 79784 142936 79812
rect 141700 79766 141752 79772
rect 141574 79716 141648 79744
rect 141344 79580 141464 79608
rect 141252 78764 141372 78792
rect 141238 78704 141294 78713
rect 141238 78639 141294 78648
rect 141252 23458 141280 78639
rect 141344 75954 141372 78764
rect 141436 78520 141464 79580
rect 141436 78492 141556 78520
rect 141424 76016 141476 76022
rect 141424 75958 141476 75964
rect 141332 75948 141384 75954
rect 141332 75890 141384 75896
rect 141332 75812 141384 75818
rect 141332 75754 141384 75760
rect 141240 23452 141292 23458
rect 141240 23394 141292 23400
rect 141344 23050 141372 75754
rect 141332 23044 141384 23050
rect 141332 22986 141384 22992
rect 140044 3052 140096 3058
rect 140044 2994 140096 3000
rect 141148 3052 141200 3058
rect 141148 2994 141200 3000
rect 140056 480 140084 2994
rect 137204 354 137232 462
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 354 141322 480
rect 141436 354 141464 75958
rect 141528 73234 141556 78492
rect 141620 76022 141648 79716
rect 141608 76016 141660 76022
rect 141608 75958 141660 75964
rect 141516 73228 141568 73234
rect 141516 73170 141568 73176
rect 141712 70394 141740 79766
rect 142172 79750 142246 79778
rect 142344 79756 142396 79762
rect 141884 79688 141936 79694
rect 141884 79630 141936 79636
rect 142068 79688 142120 79694
rect 142068 79630 142120 79636
rect 141792 79484 141844 79490
rect 141792 79426 141844 79432
rect 141804 75818 141832 79426
rect 141896 79218 141924 79630
rect 141976 79348 142028 79354
rect 141976 79290 142028 79296
rect 141884 79212 141936 79218
rect 141884 79154 141936 79160
rect 141792 75812 141844 75818
rect 141792 75754 141844 75760
rect 141988 73154 142016 79290
rect 142080 76673 142108 79630
rect 142066 76664 142122 76673
rect 142172 76634 142200 79750
rect 142344 79698 142396 79704
rect 142252 79688 142304 79694
rect 142252 79630 142304 79636
rect 142066 76599 142122 76608
rect 142160 76628 142212 76634
rect 142160 76570 142212 76576
rect 141896 73126 142016 73154
rect 141896 71806 141924 73126
rect 141884 71800 141936 71806
rect 141884 71742 141936 71748
rect 141528 70366 141740 70394
rect 141528 3330 141556 70366
rect 142160 23452 142212 23458
rect 142160 23394 142212 23400
rect 141516 3324 141568 3330
rect 141516 3266 141568 3272
rect 141210 326 141464 354
rect 142172 354 142200 23394
rect 142264 3194 142292 79630
rect 142356 76770 142384 79698
rect 142908 79694 142936 79784
rect 142988 79766 143040 79772
rect 142712 79688 142764 79694
rect 142712 79630 142764 79636
rect 142896 79688 142948 79694
rect 142896 79630 142948 79636
rect 142436 79552 142488 79558
rect 142436 79494 142488 79500
rect 142344 76764 142396 76770
rect 142344 76706 142396 76712
rect 142342 76664 142398 76673
rect 142342 76599 142398 76608
rect 142356 5234 142384 76599
rect 142344 5228 142396 5234
rect 142344 5170 142396 5176
rect 142448 5166 142476 79494
rect 142724 79336 142752 79630
rect 142896 79484 142948 79490
rect 142896 79426 142948 79432
rect 142724 79308 142844 79336
rect 142620 76628 142672 76634
rect 142620 76570 142672 76576
rect 142712 76628 142764 76634
rect 142712 76570 142764 76576
rect 142528 74996 142580 75002
rect 142528 74938 142580 74944
rect 142436 5160 142488 5166
rect 142436 5102 142488 5108
rect 142540 4894 142568 74938
rect 142632 23118 142660 76570
rect 142724 60518 142752 76570
rect 142816 67590 142844 79308
rect 142908 76634 142936 79426
rect 142896 76628 142948 76634
rect 142896 76570 142948 76576
rect 143000 75002 143028 79766
rect 143138 79744 143166 80036
rect 143092 79716 143166 79744
rect 143092 77704 143120 79716
rect 143230 79540 143258 80036
rect 143322 79642 143350 80036
rect 143414 79812 143442 80036
rect 143506 79937 143534 80036
rect 143492 79928 143548 79937
rect 143598 79898 143626 80036
rect 143690 79971 143718 80036
rect 143676 79962 143732 79971
rect 143782 79966 143810 80036
rect 143492 79863 143548 79872
rect 143586 79892 143638 79898
rect 143676 79897 143732 79906
rect 143770 79960 143822 79966
rect 143770 79902 143822 79908
rect 143586 79834 143638 79840
rect 143724 79824 143776 79830
rect 143414 79801 143488 79812
rect 143414 79792 143502 79801
rect 143414 79784 143446 79792
rect 143724 79766 143776 79772
rect 143446 79727 143502 79736
rect 143632 79756 143684 79762
rect 143632 79698 143684 79704
rect 143448 79688 143500 79694
rect 143322 79614 143396 79642
rect 143448 79630 143500 79636
rect 143540 79688 143592 79694
rect 143540 79630 143592 79636
rect 143230 79512 143304 79540
rect 143092 77676 143212 77704
rect 143184 77450 143212 77676
rect 143172 77444 143224 77450
rect 143172 77386 143224 77392
rect 143276 77353 143304 79512
rect 143368 77489 143396 79614
rect 143354 77480 143410 77489
rect 143354 77415 143410 77424
rect 143262 77344 143318 77353
rect 143262 77279 143318 77288
rect 143080 76764 143132 76770
rect 143080 76706 143132 76712
rect 142988 74996 143040 75002
rect 142988 74938 143040 74944
rect 143092 70394 143120 76706
rect 143460 73154 143488 79630
rect 143184 73126 143488 73154
rect 143552 73154 143580 79630
rect 143644 77294 143672 79698
rect 143736 77450 143764 79766
rect 143874 79744 143902 80036
rect 143966 79898 143994 80036
rect 143954 79892 144006 79898
rect 143954 79834 144006 79840
rect 144058 79744 144086 80036
rect 143828 79716 143902 79744
rect 144012 79716 144086 79744
rect 144150 79744 144178 80036
rect 144242 79937 144270 80036
rect 144228 79928 144284 79937
rect 144228 79863 144284 79872
rect 144334 79744 144362 80036
rect 144426 79898 144454 80036
rect 144518 79898 144546 80036
rect 144414 79892 144466 79898
rect 144414 79834 144466 79840
rect 144506 79892 144558 79898
rect 144506 79834 144558 79840
rect 144610 79744 144638 80036
rect 144702 79937 144730 80036
rect 144794 79966 144822 80036
rect 144886 79966 144914 80036
rect 144782 79960 144834 79966
rect 144688 79928 144744 79937
rect 144782 79902 144834 79908
rect 144874 79960 144926 79966
rect 144874 79902 144926 79908
rect 144688 79863 144744 79872
rect 144736 79824 144788 79830
rect 144828 79824 144880 79830
rect 144736 79766 144788 79772
rect 144826 79792 144828 79801
rect 144880 79792 144882 79801
rect 144150 79716 144224 79744
rect 143724 77444 143776 77450
rect 143724 77386 143776 77392
rect 143644 77266 143764 77294
rect 143552 73126 143672 73154
rect 143184 72486 143212 73126
rect 143172 72480 143224 72486
rect 143172 72422 143224 72428
rect 143092 70366 143488 70394
rect 142804 67584 142856 67590
rect 142804 67526 142856 67532
rect 142712 60512 142764 60518
rect 142712 60454 142764 60460
rect 142620 23112 142672 23118
rect 142620 23054 142672 23060
rect 142528 4888 142580 4894
rect 142528 4830 142580 4836
rect 143460 3806 143488 70366
rect 143448 3800 143500 3806
rect 143448 3742 143500 3748
rect 143644 3534 143672 73126
rect 143736 3670 143764 77266
rect 143828 76362 143856 79716
rect 143908 79620 143960 79626
rect 143908 79562 143960 79568
rect 143816 76356 143868 76362
rect 143816 76298 143868 76304
rect 143816 74724 143868 74730
rect 143816 74666 143868 74672
rect 143828 5438 143856 74666
rect 143816 5432 143868 5438
rect 143816 5374 143868 5380
rect 143920 5098 143948 79562
rect 143908 5092 143960 5098
rect 143908 5034 143960 5040
rect 144012 5030 144040 79716
rect 144092 79552 144144 79558
rect 144092 79494 144144 79500
rect 144104 77625 144132 79494
rect 144090 77616 144146 77625
rect 144090 77551 144146 77560
rect 144092 76356 144144 76362
rect 144092 76298 144144 76304
rect 144000 5024 144052 5030
rect 144000 4966 144052 4972
rect 144104 4826 144132 76298
rect 144196 74730 144224 79716
rect 144288 79716 144362 79744
rect 144564 79716 144638 79744
rect 144184 74724 144236 74730
rect 144184 74666 144236 74672
rect 144288 70394 144316 79716
rect 144368 79484 144420 79490
rect 144368 79426 144420 79432
rect 144380 78674 144408 79426
rect 144460 79212 144512 79218
rect 144460 79154 144512 79160
rect 144472 78946 144500 79154
rect 144460 78940 144512 78946
rect 144460 78882 144512 78888
rect 144368 78668 144420 78674
rect 144368 78610 144420 78616
rect 144564 77489 144592 79716
rect 144644 79620 144696 79626
rect 144644 79562 144696 79568
rect 144550 77480 144606 77489
rect 144368 77444 144420 77450
rect 144550 77415 144606 77424
rect 144368 77386 144420 77392
rect 144380 73154 144408 77386
rect 144550 76664 144606 76673
rect 144550 76599 144606 76608
rect 144380 73126 144500 73154
rect 144196 70366 144316 70394
rect 144196 58818 144224 70366
rect 144184 58812 144236 58818
rect 144184 58754 144236 58760
rect 144092 4820 144144 4826
rect 144092 4762 144144 4768
rect 144472 3874 144500 73126
rect 144460 3868 144512 3874
rect 144460 3810 144512 3816
rect 143724 3664 143776 3670
rect 143724 3606 143776 3612
rect 143632 3528 143684 3534
rect 143632 3470 143684 3476
rect 144564 3466 144592 76599
rect 144656 75682 144684 79562
rect 144644 75676 144696 75682
rect 144644 75618 144696 75624
rect 144748 71262 144776 79766
rect 144826 79727 144882 79736
rect 144978 79676 145006 80036
rect 145070 79830 145098 80036
rect 145058 79824 145110 79830
rect 145058 79766 145110 79772
rect 145162 79676 145190 80036
rect 145254 79966 145282 80036
rect 145242 79960 145294 79966
rect 145242 79902 145294 79908
rect 144840 79648 145006 79676
rect 145116 79648 145190 79676
rect 145346 79676 145374 80036
rect 145438 79744 145466 80036
rect 145530 79966 145558 80036
rect 145518 79960 145570 79966
rect 145518 79902 145570 79908
rect 145438 79716 145512 79744
rect 145346 79648 145420 79676
rect 144840 77246 144868 79648
rect 145116 79506 145144 79648
rect 145024 79478 145144 79506
rect 145288 79552 145340 79558
rect 145288 79494 145340 79500
rect 145196 79484 145248 79490
rect 144920 79416 144972 79422
rect 144920 79358 144972 79364
rect 144932 78946 144960 79358
rect 144920 78940 144972 78946
rect 144920 78882 144972 78888
rect 144918 77480 144974 77489
rect 144918 77415 144974 77424
rect 144828 77240 144880 77246
rect 144828 77182 144880 77188
rect 144736 71256 144788 71262
rect 144736 71198 144788 71204
rect 144932 6118 144960 77415
rect 145024 26110 145052 79478
rect 145196 79426 145248 79432
rect 145104 79416 145156 79422
rect 145104 79358 145156 79364
rect 145116 77294 145144 79358
rect 145208 78062 145236 79426
rect 145196 78056 145248 78062
rect 145196 77998 145248 78004
rect 145116 77266 145236 77294
rect 145104 77172 145156 77178
rect 145104 77114 145156 77120
rect 145116 26994 145144 77114
rect 145208 32638 145236 77266
rect 145300 32706 145328 79494
rect 145392 77994 145420 79648
rect 145484 78130 145512 79716
rect 145622 79676 145650 80036
rect 145714 79744 145742 80036
rect 145806 79812 145834 80036
rect 145898 79937 145926 80036
rect 145884 79928 145940 79937
rect 145884 79863 145940 79872
rect 145806 79784 145880 79812
rect 145714 79716 145788 79744
rect 145576 79648 145650 79676
rect 145472 78124 145524 78130
rect 145472 78066 145524 78072
rect 145380 77988 145432 77994
rect 145380 77930 145432 77936
rect 145380 76968 145432 76974
rect 145380 76910 145432 76916
rect 145288 32700 145340 32706
rect 145288 32642 145340 32648
rect 145196 32632 145248 32638
rect 145196 32574 145248 32580
rect 145392 32570 145420 76910
rect 145472 76424 145524 76430
rect 145472 76366 145524 76372
rect 145484 62830 145512 76366
rect 145576 68882 145604 79648
rect 145656 79552 145708 79558
rect 145656 79494 145708 79500
rect 145668 77489 145696 79494
rect 145654 77480 145710 77489
rect 145654 77415 145710 77424
rect 145760 77178 145788 79716
rect 145852 79422 145880 79784
rect 145990 79608 146018 80036
rect 146082 79676 146110 80036
rect 146174 79898 146202 80036
rect 146266 79898 146294 80036
rect 146358 79898 146386 80036
rect 146162 79892 146214 79898
rect 146162 79834 146214 79840
rect 146254 79892 146306 79898
rect 146254 79834 146306 79840
rect 146346 79892 146398 79898
rect 146346 79834 146398 79840
rect 146450 79778 146478 80036
rect 146542 79801 146570 80036
rect 146634 79898 146662 80036
rect 146622 79892 146674 79898
rect 146622 79834 146674 79840
rect 146404 79750 146478 79778
rect 146528 79792 146584 79801
rect 146208 79688 146260 79694
rect 146082 79648 146156 79676
rect 145990 79580 146064 79608
rect 145932 79484 145984 79490
rect 145932 79426 145984 79432
rect 145840 79416 145892 79422
rect 145840 79358 145892 79364
rect 145748 77172 145800 77178
rect 145748 77114 145800 77120
rect 145944 75818 145972 79426
rect 146036 76430 146064 79580
rect 146128 76974 146156 79648
rect 146208 79630 146260 79636
rect 146220 77489 146248 79630
rect 146300 79484 146352 79490
rect 146300 79426 146352 79432
rect 146206 77480 146262 77489
rect 146206 77415 146262 77424
rect 146208 77172 146260 77178
rect 146208 77114 146260 77120
rect 146116 76968 146168 76974
rect 146116 76910 146168 76916
rect 146024 76424 146076 76430
rect 146024 76366 146076 76372
rect 145932 75812 145984 75818
rect 145932 75754 145984 75760
rect 145564 68876 145616 68882
rect 145564 68818 145616 68824
rect 145564 67584 145616 67590
rect 145564 67526 145616 67532
rect 145472 62824 145524 62830
rect 145472 62766 145524 62772
rect 145380 32564 145432 32570
rect 145380 32506 145432 32512
rect 145104 26988 145156 26994
rect 145104 26930 145156 26936
rect 145012 26104 145064 26110
rect 145012 26046 145064 26052
rect 145012 23044 145064 23050
rect 145012 22986 145064 22992
rect 145024 16574 145052 22986
rect 145024 16546 145512 16574
rect 144920 6112 144972 6118
rect 144920 6054 144972 6060
rect 144736 4140 144788 4146
rect 144736 4082 144788 4088
rect 144552 3460 144604 3466
rect 144552 3402 144604 3408
rect 143540 3324 143592 3330
rect 143540 3266 143592 3272
rect 142252 3188 142304 3194
rect 142252 3130 142304 3136
rect 143552 480 143580 3266
rect 144748 480 144776 4082
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 141210 -960 141322 326
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 145576 3058 145604 67526
rect 146220 18698 146248 77114
rect 146208 18692 146260 18698
rect 146208 18634 146260 18640
rect 146312 9178 146340 79426
rect 146404 76294 146432 79750
rect 146726 79778 146754 80036
rect 146818 79898 146846 80036
rect 146806 79892 146858 79898
rect 146806 79834 146858 79840
rect 146528 79727 146584 79736
rect 146680 79750 146754 79778
rect 146910 79778 146938 80036
rect 147002 79966 147030 80036
rect 146990 79960 147042 79966
rect 147094 79937 147122 80036
rect 147186 79966 147214 80036
rect 147174 79960 147226 79966
rect 146990 79902 147042 79908
rect 147080 79928 147136 79937
rect 147174 79902 147226 79908
rect 147278 79898 147306 80036
rect 147370 79898 147398 80036
rect 147462 79971 147490 80036
rect 147448 79962 147504 79971
rect 147080 79863 147136 79872
rect 147266 79892 147318 79898
rect 147266 79834 147318 79840
rect 147358 79892 147410 79898
rect 147448 79897 147504 79906
rect 147358 79834 147410 79840
rect 147554 79830 147582 80036
rect 147542 79824 147594 79830
rect 146910 79750 147076 79778
rect 147542 79766 147594 79772
rect 146680 79472 146708 79750
rect 146944 79688 146996 79694
rect 146864 79648 146944 79676
rect 146760 79552 146812 79558
rect 146760 79494 146812 79500
rect 146588 79444 146708 79472
rect 146484 79416 146536 79422
rect 146484 79358 146536 79364
rect 146392 76288 146444 76294
rect 146392 76230 146444 76236
rect 146392 76152 146444 76158
rect 146392 76094 146444 76100
rect 146404 12442 146432 76094
rect 146496 23390 146524 79358
rect 146588 78538 146616 79444
rect 146576 78532 146628 78538
rect 146576 78474 146628 78480
rect 146574 77344 146630 77353
rect 146574 77279 146630 77288
rect 146484 23384 146536 23390
rect 146484 23326 146536 23332
rect 146588 23322 146616 77279
rect 146666 76664 146722 76673
rect 146666 76599 146722 76608
rect 146680 23458 146708 76599
rect 146772 28082 146800 79494
rect 146864 28150 146892 79648
rect 146944 79630 146996 79636
rect 147048 74534 147076 79750
rect 147404 79756 147456 79762
rect 147404 79698 147456 79704
rect 147220 79688 147272 79694
rect 147220 79630 147272 79636
rect 147128 79620 147180 79626
rect 147128 79562 147180 79568
rect 147140 76566 147168 79562
rect 147128 76560 147180 76566
rect 147128 76502 147180 76508
rect 147232 76158 147260 79630
rect 147312 78124 147364 78130
rect 147312 78066 147364 78072
rect 147220 76152 147272 76158
rect 147220 76094 147272 76100
rect 147324 74534 147352 78066
rect 147416 77353 147444 79698
rect 147496 79688 147548 79694
rect 147646 79676 147674 80036
rect 147738 79830 147766 80036
rect 147830 79898 147858 80036
rect 147922 79966 147950 80036
rect 147910 79960 147962 79966
rect 147910 79902 147962 79908
rect 147818 79892 147870 79898
rect 147818 79834 147870 79840
rect 147726 79824 147778 79830
rect 147726 79766 147778 79772
rect 148014 79744 148042 80036
rect 148106 79812 148134 80036
rect 148198 79966 148226 80036
rect 148290 79966 148318 80036
rect 148382 79966 148410 80036
rect 148474 79971 148502 80036
rect 148186 79960 148238 79966
rect 148186 79902 148238 79908
rect 148278 79960 148330 79966
rect 148278 79902 148330 79908
rect 148370 79960 148422 79966
rect 148370 79902 148422 79908
rect 148460 79962 148516 79971
rect 148460 79897 148516 79906
rect 148566 79898 148594 80036
rect 148658 79971 148686 80036
rect 148644 79962 148700 79971
rect 148750 79966 148778 80036
rect 148554 79892 148606 79898
rect 148644 79897 148700 79906
rect 148738 79960 148790 79966
rect 148842 79937 148870 80036
rect 148738 79902 148790 79908
rect 148828 79928 148884 79937
rect 148934 79898 148962 80036
rect 149026 79898 149054 80036
rect 149118 79971 149146 80036
rect 149104 79962 149160 79971
rect 148828 79863 148884 79872
rect 148922 79892 148974 79898
rect 148554 79834 148606 79840
rect 148922 79834 148974 79840
rect 149014 79892 149066 79898
rect 149104 79897 149160 79906
rect 149210 79898 149238 80036
rect 149014 79834 149066 79840
rect 149198 79892 149250 79898
rect 149198 79834 149250 79840
rect 148784 79824 148836 79830
rect 148106 79784 148180 79812
rect 148014 79716 148088 79744
rect 147772 79688 147824 79694
rect 147646 79648 147720 79676
rect 147496 79630 147548 79636
rect 147508 77489 147536 79630
rect 147588 77988 147640 77994
rect 147588 77930 147640 77936
rect 147494 77480 147550 77489
rect 147494 77415 147550 77424
rect 147402 77344 147458 77353
rect 147402 77279 147458 77288
rect 146956 74506 147076 74534
rect 147140 74506 147352 74534
rect 146956 28218 146984 74506
rect 147140 70394 147168 74506
rect 147600 70394 147628 77930
rect 147692 77178 147720 79648
rect 147772 79630 147824 79636
rect 147784 77294 147812 79630
rect 148060 77654 148088 79716
rect 148048 77648 148100 77654
rect 148048 77590 148100 77596
rect 147956 77580 148008 77586
rect 147956 77522 148008 77528
rect 147784 77266 147904 77294
rect 147680 77172 147732 77178
rect 147680 77114 147732 77120
rect 147772 77172 147824 77178
rect 147772 77114 147824 77120
rect 147680 76628 147732 76634
rect 147680 76570 147732 76576
rect 147048 70366 147168 70394
rect 147232 70366 147628 70394
rect 146944 28212 146996 28218
rect 146944 28154 146996 28160
rect 146852 28144 146904 28150
rect 146852 28086 146904 28092
rect 146760 28076 146812 28082
rect 146760 28018 146812 28024
rect 146668 23452 146720 23458
rect 146668 23394 146720 23400
rect 146576 23316 146628 23322
rect 146576 23258 146628 23264
rect 147048 14278 147076 70366
rect 147036 14272 147088 14278
rect 147036 14214 147088 14220
rect 146392 12436 146444 12442
rect 146392 12378 146444 12384
rect 146300 9172 146352 9178
rect 146300 9114 146352 9120
rect 147128 3596 147180 3602
rect 147128 3538 147180 3544
rect 145564 3052 145616 3058
rect 145564 2994 145616 3000
rect 147140 480 147168 3538
rect 147232 3262 147260 70366
rect 147692 3398 147720 76570
rect 147784 4078 147812 77114
rect 147876 4962 147904 77266
rect 147968 12306 147996 77522
rect 148152 77432 148180 79784
rect 149302 79812 149330 80036
rect 149394 79966 149422 80036
rect 149382 79960 149434 79966
rect 149382 79902 149434 79908
rect 149486 79812 149514 80036
rect 149578 79971 149606 80036
rect 149564 79962 149620 79971
rect 149564 79897 149620 79906
rect 149670 79898 149698 80036
rect 149762 79937 149790 80036
rect 149748 79928 149804 79937
rect 149658 79892 149710 79898
rect 149748 79863 149804 79872
rect 149658 79834 149710 79840
rect 148784 79766 148836 79772
rect 149058 79792 149114 79801
rect 148324 79756 148376 79762
rect 148324 79698 148376 79704
rect 148232 79688 148284 79694
rect 148232 79630 148284 79636
rect 148244 77586 148272 79630
rect 148232 77580 148284 77586
rect 148232 77522 148284 77528
rect 148060 77404 148180 77432
rect 148060 77178 148088 77404
rect 148048 77172 148100 77178
rect 148048 77114 148100 77120
rect 148046 76664 148102 76673
rect 148336 76616 148364 79698
rect 148416 79688 148468 79694
rect 148468 79648 148548 79676
rect 148416 79630 148468 79636
rect 148416 77648 148468 77654
rect 148416 77590 148468 77596
rect 148046 76599 148102 76608
rect 147956 12300 148008 12306
rect 147956 12242 148008 12248
rect 148060 12238 148088 76599
rect 148244 76588 148364 76616
rect 148140 76560 148192 76566
rect 148140 76502 148192 76508
rect 148152 12374 148180 76502
rect 148244 17678 148272 76588
rect 148428 73154 148456 77590
rect 148520 76634 148548 79648
rect 148600 79620 148652 79626
rect 148600 79562 148652 79568
rect 148692 79620 148744 79626
rect 148692 79562 148744 79568
rect 148508 76628 148560 76634
rect 148508 76570 148560 76576
rect 148612 74526 148640 79562
rect 148704 77586 148732 79562
rect 148692 77580 148744 77586
rect 148692 77522 148744 77528
rect 148796 76129 148824 79766
rect 148876 79756 148928 79762
rect 149302 79784 149376 79812
rect 149486 79784 149560 79812
rect 149058 79727 149114 79736
rect 149152 79756 149204 79762
rect 148876 79698 148928 79704
rect 148782 76120 148838 76129
rect 148782 76055 148838 76064
rect 148888 75993 148916 79698
rect 148968 79416 149020 79422
rect 148968 79358 149020 79364
rect 148874 75984 148930 75993
rect 148874 75919 148930 75928
rect 148980 75750 149008 79358
rect 149072 75954 149100 79727
rect 149152 79698 149204 79704
rect 149060 75948 149112 75954
rect 149060 75890 149112 75896
rect 148968 75744 149020 75750
rect 148968 75686 149020 75692
rect 148600 74520 148652 74526
rect 148600 74462 148652 74468
rect 148336 73126 148456 73154
rect 148336 60246 148364 73126
rect 148416 60512 148468 60518
rect 148416 60454 148468 60460
rect 148324 60240 148376 60246
rect 148324 60182 148376 60188
rect 148232 17672 148284 17678
rect 148232 17614 148284 17620
rect 148140 12368 148192 12374
rect 148140 12310 148192 12316
rect 148048 12232 148100 12238
rect 148048 12174 148100 12180
rect 147864 4956 147916 4962
rect 147864 4898 147916 4904
rect 148428 4146 148456 60454
rect 149060 23112 149112 23118
rect 149060 23054 149112 23060
rect 148416 4140 148468 4146
rect 148416 4082 148468 4088
rect 147772 4072 147824 4078
rect 147772 4014 147824 4020
rect 148322 3632 148378 3641
rect 148322 3567 148378 3576
rect 147680 3392 147732 3398
rect 147680 3334 147732 3340
rect 147220 3256 147272 3262
rect 147220 3198 147272 3204
rect 148336 480 148364 3567
rect 149072 3482 149100 23054
rect 149164 4010 149192 79698
rect 149348 79676 149376 79784
rect 149256 79648 149376 79676
rect 149428 79688 149480 79694
rect 149256 79490 149284 79648
rect 149532 79676 149560 79784
rect 149854 79778 149882 80036
rect 149946 79966 149974 80036
rect 150038 79966 150066 80036
rect 149934 79960 149986 79966
rect 149934 79902 149986 79908
rect 150026 79960 150078 79966
rect 150026 79902 150078 79908
rect 149808 79750 149882 79778
rect 149980 79756 150032 79762
rect 149532 79648 149652 79676
rect 149428 79630 149480 79636
rect 149244 79484 149296 79490
rect 149244 79426 149296 79432
rect 149336 79416 149388 79422
rect 149336 79358 149388 79364
rect 149244 79348 149296 79354
rect 149244 79290 149296 79296
rect 149256 79121 149284 79290
rect 149242 79112 149298 79121
rect 149242 79047 149298 79056
rect 149244 75948 149296 75954
rect 149244 75890 149296 75896
rect 149256 6798 149284 75890
rect 149348 9110 149376 79358
rect 149440 76809 149468 79630
rect 149520 79484 149572 79490
rect 149520 79426 149572 79432
rect 149426 76800 149482 76809
rect 149426 76735 149482 76744
rect 149426 76120 149482 76129
rect 149426 76055 149482 76064
rect 149440 12102 149468 76055
rect 149532 12170 149560 79426
rect 149624 76566 149652 79648
rect 149808 79422 149836 79750
rect 150130 79744 150158 80036
rect 150222 79898 150250 80036
rect 150314 79971 150342 80036
rect 150300 79962 150356 79971
rect 150210 79892 150262 79898
rect 150300 79897 150356 79906
rect 150406 79898 150434 80036
rect 150498 79898 150526 80036
rect 150210 79834 150262 79840
rect 150394 79892 150446 79898
rect 150394 79834 150446 79840
rect 150486 79892 150538 79898
rect 150486 79834 150538 79840
rect 150590 79830 150618 80036
rect 150682 79898 150710 80036
rect 150774 79971 150802 80036
rect 150760 79962 150816 79971
rect 150670 79892 150722 79898
rect 150760 79897 150816 79906
rect 150670 79834 150722 79840
rect 150578 79824 150630 79830
rect 150578 79766 150630 79772
rect 149980 79698 150032 79704
rect 150084 79716 150158 79744
rect 150716 79756 150768 79762
rect 149888 79688 149940 79694
rect 149888 79630 149940 79636
rect 149796 79416 149848 79422
rect 149796 79358 149848 79364
rect 149612 76560 149664 76566
rect 149612 76502 149664 76508
rect 149900 76430 149928 79630
rect 149612 76424 149664 76430
rect 149612 76366 149664 76372
rect 149888 76424 149940 76430
rect 149888 76366 149940 76372
rect 149624 15978 149652 76366
rect 149888 76288 149940 76294
rect 149888 76230 149940 76236
rect 149702 75984 149758 75993
rect 149702 75919 149758 75928
rect 149716 19922 149744 75919
rect 149900 70394 149928 76230
rect 149992 75993 150020 79698
rect 150084 76673 150112 79716
rect 150866 79744 150894 80036
rect 150958 79971 150986 80036
rect 150944 79962 151000 79971
rect 150944 79897 151000 79906
rect 151050 79898 151078 80036
rect 151142 79966 151170 80036
rect 151130 79960 151182 79966
rect 151130 79902 151182 79908
rect 151234 79898 151262 80036
rect 151326 79966 151354 80036
rect 151418 79966 151446 80036
rect 151510 79966 151538 80036
rect 151314 79960 151366 79966
rect 151314 79902 151366 79908
rect 151406 79960 151458 79966
rect 151406 79902 151458 79908
rect 151498 79960 151550 79966
rect 151498 79902 151550 79908
rect 151038 79892 151090 79898
rect 151038 79834 151090 79840
rect 151222 79892 151274 79898
rect 151222 79834 151274 79840
rect 151602 79778 151630 80036
rect 151694 79971 151722 80036
rect 151680 79962 151736 79971
rect 151680 79897 151736 79906
rect 151786 79898 151814 80036
rect 151878 79898 151906 80036
rect 151970 79966 151998 80036
rect 151958 79960 152010 79966
rect 151958 79902 152010 79908
rect 151774 79892 151826 79898
rect 151774 79834 151826 79840
rect 151866 79892 151918 79898
rect 151866 79834 151918 79840
rect 150716 79698 150768 79704
rect 150820 79716 150894 79744
rect 151084 79756 151136 79762
rect 150256 79688 150308 79694
rect 150256 79630 150308 79636
rect 150624 79688 150676 79694
rect 150624 79630 150676 79636
rect 150164 79552 150216 79558
rect 150164 79494 150216 79500
rect 150070 76664 150126 76673
rect 150070 76599 150126 76608
rect 150072 76560 150124 76566
rect 150072 76502 150124 76508
rect 149978 75984 150034 75993
rect 149978 75919 150034 75928
rect 149900 70366 150020 70394
rect 149704 19916 149756 19922
rect 149704 19858 149756 19864
rect 149612 15972 149664 15978
rect 149612 15914 149664 15920
rect 149520 12164 149572 12170
rect 149520 12106 149572 12112
rect 149428 12096 149480 12102
rect 149428 12038 149480 12044
rect 149336 9104 149388 9110
rect 149336 9046 149388 9052
rect 149992 6866 150020 70366
rect 149980 6860 150032 6866
rect 149980 6802 150032 6808
rect 149244 6792 149296 6798
rect 149244 6734 149296 6740
rect 149244 5432 149296 5438
rect 149244 5374 149296 5380
rect 149152 4004 149204 4010
rect 149152 3946 149204 3952
rect 149256 3602 149284 5374
rect 150084 3777 150112 76502
rect 150176 74322 150204 79494
rect 150164 74316 150216 74322
rect 150164 74258 150216 74264
rect 150268 74089 150296 79630
rect 150440 79552 150492 79558
rect 150440 79494 150492 79500
rect 150254 74080 150310 74089
rect 150254 74015 150310 74024
rect 150452 3942 150480 79494
rect 150636 77194 150664 79630
rect 150728 78606 150756 79698
rect 150716 78600 150768 78606
rect 150716 78542 150768 78548
rect 150820 78130 150848 79716
rect 151084 79698 151136 79704
rect 151176 79756 151228 79762
rect 151176 79698 151228 79704
rect 151268 79756 151320 79762
rect 151268 79698 151320 79704
rect 151556 79750 151630 79778
rect 150900 79620 150952 79626
rect 150900 79562 150952 79568
rect 150808 78124 150860 78130
rect 150808 78066 150860 78072
rect 150636 77166 150848 77194
rect 150624 77036 150676 77042
rect 150624 76978 150676 76984
rect 150636 76106 150664 76978
rect 150544 76078 150664 76106
rect 150820 76106 150848 77166
rect 150912 77042 150940 79562
rect 150990 78296 151046 78305
rect 150990 78231 151046 78240
rect 150900 77036 150952 77042
rect 150900 76978 150952 76984
rect 150820 76078 150940 76106
rect 150440 3936 150492 3942
rect 150440 3878 150492 3884
rect 150070 3768 150126 3777
rect 150070 3703 150126 3712
rect 150544 3641 150572 76078
rect 150624 76016 150676 76022
rect 150624 75958 150676 75964
rect 150714 75984 150770 75993
rect 150636 6730 150664 75958
rect 150714 75919 150770 75928
rect 150808 75948 150860 75954
rect 150728 14346 150756 75919
rect 150808 75890 150860 75896
rect 150820 14414 150848 75890
rect 150912 20670 150940 76078
rect 150900 20664 150952 20670
rect 150900 20606 150952 20612
rect 151004 20602 151032 78231
rect 150992 20596 151044 20602
rect 150992 20538 151044 20544
rect 151096 20534 151124 79698
rect 151188 75954 151216 79698
rect 151280 78169 151308 79698
rect 151360 79688 151412 79694
rect 151360 79630 151412 79636
rect 151266 78160 151322 78169
rect 151266 78095 151322 78104
rect 151372 76022 151400 79630
rect 151452 79620 151504 79626
rect 151452 79562 151504 79568
rect 151464 76906 151492 79562
rect 151452 76900 151504 76906
rect 151452 76842 151504 76848
rect 151360 76016 151412 76022
rect 151360 75958 151412 75964
rect 151176 75948 151228 75954
rect 151176 75890 151228 75896
rect 151556 70394 151584 79750
rect 151728 79688 151780 79694
rect 151728 79630 151780 79636
rect 151912 79688 151964 79694
rect 152062 79676 152090 80036
rect 152154 79830 152182 80036
rect 152246 79898 152274 80036
rect 152338 79971 152366 80036
rect 152324 79962 152380 79971
rect 152234 79892 152286 79898
rect 152324 79897 152380 79906
rect 152430 79898 152458 80036
rect 152522 79966 152550 80036
rect 152614 79966 152642 80036
rect 152510 79960 152562 79966
rect 152510 79902 152562 79908
rect 152602 79960 152654 79966
rect 152706 79937 152734 80036
rect 152798 79966 152826 80036
rect 152890 79971 152918 80036
rect 152786 79960 152838 79966
rect 152602 79902 152654 79908
rect 152692 79928 152748 79937
rect 152234 79834 152286 79840
rect 152418 79892 152470 79898
rect 152786 79902 152838 79908
rect 152876 79962 152932 79971
rect 152982 79966 153010 80036
rect 153074 79966 153102 80036
rect 153166 79966 153194 80036
rect 153258 79966 153286 80036
rect 152876 79897 152932 79906
rect 152970 79960 153022 79966
rect 152970 79902 153022 79908
rect 153062 79960 153114 79966
rect 153062 79902 153114 79908
rect 153154 79960 153206 79966
rect 153154 79902 153206 79908
rect 153246 79960 153298 79966
rect 153246 79902 153298 79908
rect 152692 79863 152748 79872
rect 152418 79834 152470 79840
rect 152142 79824 152194 79830
rect 153350 79812 153378 80036
rect 153442 79971 153470 80036
rect 153428 79962 153484 79971
rect 153428 79897 153484 79906
rect 153534 79830 153562 80036
rect 153626 79830 153654 80036
rect 153718 79937 153746 80036
rect 153704 79928 153760 79937
rect 153704 79863 153760 79872
rect 153522 79824 153574 79830
rect 153350 79784 153424 79812
rect 152142 79766 152194 79772
rect 152280 79756 152332 79762
rect 152280 79698 152332 79704
rect 152372 79756 152424 79762
rect 152372 79698 152424 79704
rect 152648 79756 152700 79762
rect 152648 79698 152700 79704
rect 152832 79756 152884 79762
rect 152832 79698 152884 79704
rect 153108 79756 153160 79762
rect 153108 79698 153160 79704
rect 151912 79630 151964 79636
rect 152016 79648 152090 79676
rect 151636 79620 151688 79626
rect 151636 79562 151688 79568
rect 151648 75993 151676 79562
rect 151634 75984 151690 75993
rect 151740 75954 151768 79630
rect 151820 79620 151872 79626
rect 151820 79562 151872 79568
rect 151634 75919 151690 75928
rect 151728 75948 151780 75954
rect 151728 75890 151780 75896
rect 151188 70366 151584 70394
rect 151084 20528 151136 20534
rect 151084 20470 151136 20476
rect 151188 20466 151216 70366
rect 151176 20460 151228 20466
rect 151176 20402 151228 20408
rect 150808 14408 150860 14414
rect 150808 14350 150860 14356
rect 150716 14340 150768 14346
rect 150716 14282 150768 14288
rect 150624 6724 150676 6730
rect 150624 6666 150676 6672
rect 151832 6662 151860 79562
rect 151924 75546 151952 79630
rect 152016 79540 152044 79648
rect 152188 79552 152240 79558
rect 152016 79512 152136 79540
rect 152004 76016 152056 76022
rect 152004 75958 152056 75964
rect 151912 75540 151964 75546
rect 151912 75482 151964 75488
rect 151912 74044 151964 74050
rect 151912 73986 151964 73992
rect 151820 6656 151872 6662
rect 151820 6598 151872 6604
rect 151924 6594 151952 73986
rect 152016 15026 152044 75958
rect 152108 15162 152136 79512
rect 152188 79494 152240 79500
rect 152200 77217 152228 79494
rect 152186 77208 152242 77217
rect 152186 77143 152242 77152
rect 152186 75984 152242 75993
rect 152186 75919 152242 75928
rect 152096 15156 152148 15162
rect 152096 15098 152148 15104
rect 152200 15094 152228 75919
rect 152292 20398 152320 79698
rect 152384 23186 152412 79698
rect 152556 79620 152608 79626
rect 152556 79562 152608 79568
rect 152464 75948 152516 75954
rect 152464 75890 152516 75896
rect 152476 23254 152504 75890
rect 152568 74050 152596 79562
rect 152660 79506 152688 79698
rect 152660 79478 152780 79506
rect 152648 79416 152700 79422
rect 152648 79358 152700 79364
rect 152556 74044 152608 74050
rect 152556 73986 152608 73992
rect 152660 70394 152688 79358
rect 152752 76022 152780 79478
rect 152740 76016 152792 76022
rect 152844 75993 152872 79698
rect 153016 79484 153068 79490
rect 153016 79426 153068 79432
rect 153028 76022 153056 79426
rect 153120 76129 153148 79698
rect 153292 79688 153344 79694
rect 153292 79630 153344 79636
rect 153200 79552 153252 79558
rect 153200 79494 153252 79500
rect 153106 76120 153162 76129
rect 153106 76055 153162 76064
rect 153016 76016 153068 76022
rect 152740 75958 152792 75964
rect 152830 75984 152886 75993
rect 153016 75958 153068 75964
rect 153212 75954 153240 79494
rect 153304 76974 153332 79630
rect 153396 78928 153424 79784
rect 153522 79766 153574 79772
rect 153614 79824 153666 79830
rect 153810 79812 153838 80036
rect 153902 79966 153930 80036
rect 153994 79966 154022 80036
rect 154086 79966 154114 80036
rect 154178 79966 154206 80036
rect 154270 79966 154298 80036
rect 154362 79966 154390 80036
rect 154454 79971 154482 80036
rect 153890 79960 153942 79966
rect 153890 79902 153942 79908
rect 153982 79960 154034 79966
rect 153982 79902 154034 79908
rect 154074 79960 154126 79966
rect 154074 79902 154126 79908
rect 154166 79960 154218 79966
rect 154166 79902 154218 79908
rect 154258 79960 154310 79966
rect 154258 79902 154310 79908
rect 154350 79960 154402 79966
rect 154350 79902 154402 79908
rect 154440 79962 154496 79971
rect 154546 79966 154574 80036
rect 154638 79966 154666 80036
rect 154730 79966 154758 80036
rect 154440 79897 154496 79906
rect 154534 79960 154586 79966
rect 154534 79902 154586 79908
rect 154626 79960 154678 79966
rect 154626 79902 154678 79908
rect 154718 79960 154770 79966
rect 154718 79902 154770 79908
rect 153764 79784 153838 79812
rect 154822 79812 154850 80036
rect 154914 79937 154942 80036
rect 155006 79966 155034 80036
rect 155098 79966 155126 80036
rect 155190 79966 155218 80036
rect 155282 79966 155310 80036
rect 155374 79971 155402 80036
rect 154994 79960 155046 79966
rect 154900 79928 154956 79937
rect 154994 79902 155046 79908
rect 155086 79960 155138 79966
rect 155086 79902 155138 79908
rect 155178 79960 155230 79966
rect 155178 79902 155230 79908
rect 155270 79960 155322 79966
rect 155270 79902 155322 79908
rect 155360 79962 155416 79971
rect 155466 79966 155494 80036
rect 155558 79971 155586 80036
rect 155360 79897 155416 79906
rect 155454 79960 155506 79966
rect 155454 79902 155506 79908
rect 155544 79962 155600 79971
rect 155544 79897 155600 79906
rect 154900 79863 154956 79872
rect 155132 79824 155184 79830
rect 154822 79784 154896 79812
rect 153764 79778 153792 79784
rect 153614 79766 153666 79772
rect 153718 79750 153792 79778
rect 154028 79756 154080 79762
rect 153568 79688 153620 79694
rect 153718 79676 153746 79750
rect 154028 79698 154080 79704
rect 154304 79756 154356 79762
rect 154304 79698 154356 79704
rect 154396 79756 154448 79762
rect 154396 79698 154448 79704
rect 154672 79756 154724 79762
rect 154672 79698 154724 79704
rect 153568 79630 153620 79636
rect 153672 79648 153746 79676
rect 153844 79688 153896 79694
rect 153396 78900 153516 78928
rect 153292 76968 153344 76974
rect 153292 76910 153344 76916
rect 153384 76288 153436 76294
rect 153384 76230 153436 76236
rect 153292 76220 153344 76226
rect 153292 76162 153344 76168
rect 152830 75919 152886 75928
rect 153200 75948 153252 75954
rect 153200 75890 153252 75896
rect 153200 75608 153252 75614
rect 153200 75550 153252 75556
rect 152660 70366 152780 70394
rect 152752 26042 152780 70366
rect 152740 26036 152792 26042
rect 152740 25978 152792 25984
rect 152464 23248 152516 23254
rect 152464 23190 152516 23196
rect 152372 23180 152424 23186
rect 152372 23122 152424 23128
rect 152280 20392 152332 20398
rect 152280 20334 152332 20340
rect 152188 15088 152240 15094
rect 152188 15030 152240 15036
rect 152004 15020 152056 15026
rect 152004 14962 152056 14968
rect 151912 6588 151964 6594
rect 151912 6530 151964 6536
rect 153212 6322 153240 75550
rect 153304 6390 153332 76162
rect 153396 6458 153424 76230
rect 153488 6526 153516 78900
rect 153580 76294 153608 79630
rect 153568 76288 153620 76294
rect 153568 76230 153620 76236
rect 153566 75984 153622 75993
rect 153566 75919 153622 75928
rect 153580 14958 153608 75919
rect 153672 20330 153700 79648
rect 153844 79630 153896 79636
rect 153752 79552 153804 79558
rect 153752 79494 153804 79500
rect 153764 77081 153792 79494
rect 153750 77072 153806 77081
rect 153750 77007 153806 77016
rect 153752 76968 153804 76974
rect 153752 76910 153804 76916
rect 153764 23118 153792 76910
rect 153856 76226 153884 79630
rect 153936 79620 153988 79626
rect 153936 79562 153988 79568
rect 153844 76220 153896 76226
rect 153844 76162 153896 76168
rect 153948 76106 153976 79562
rect 153856 76078 153976 76106
rect 153752 23112 153804 23118
rect 153752 23054 153804 23060
rect 153856 22982 153884 76078
rect 153936 76016 153988 76022
rect 153936 75958 153988 75964
rect 153948 23050 153976 75958
rect 154040 75614 154068 79698
rect 154212 79484 154264 79490
rect 154212 79426 154264 79432
rect 154224 78878 154252 79426
rect 154212 78872 154264 78878
rect 154212 78814 154264 78820
rect 154316 77081 154344 79698
rect 154408 77761 154436 79698
rect 154488 79688 154540 79694
rect 154488 79630 154540 79636
rect 154394 77752 154450 77761
rect 154394 77687 154450 77696
rect 154302 77072 154358 77081
rect 154302 77007 154358 77016
rect 154500 75993 154528 79630
rect 154580 79620 154632 79626
rect 154580 79562 154632 79568
rect 154592 78470 154620 79562
rect 154580 78464 154632 78470
rect 154580 78406 154632 78412
rect 154486 75984 154542 75993
rect 154212 75948 154264 75954
rect 154486 75919 154542 75928
rect 154212 75890 154264 75896
rect 154028 75608 154080 75614
rect 154028 75550 154080 75556
rect 154224 64874 154252 75890
rect 154684 74186 154712 79698
rect 154672 74180 154724 74186
rect 154672 74122 154724 74128
rect 154868 71774 154896 79784
rect 155132 79766 155184 79772
rect 155314 79792 155370 79801
rect 154948 79756 155000 79762
rect 154948 79698 155000 79704
rect 154776 71746 154896 71774
rect 154776 71602 154804 71746
rect 154764 71596 154816 71602
rect 154764 71538 154816 71544
rect 154960 70394 154988 79698
rect 155040 79620 155092 79626
rect 155040 79562 155092 79568
rect 155052 75954 155080 79562
rect 155040 75948 155092 75954
rect 155040 75890 155092 75896
rect 155144 71774 155172 79766
rect 155650 79778 155678 80036
rect 155742 79898 155770 80036
rect 155834 79971 155862 80036
rect 155820 79962 155876 79971
rect 155730 79892 155782 79898
rect 155820 79897 155876 79906
rect 155926 79898 155954 80036
rect 156018 79898 156046 80036
rect 156110 79966 156138 80036
rect 156202 79966 156230 80036
rect 156294 79966 156322 80036
rect 156098 79960 156150 79966
rect 156098 79902 156150 79908
rect 156190 79960 156242 79966
rect 156190 79902 156242 79908
rect 156282 79960 156334 79966
rect 156282 79902 156334 79908
rect 156386 79898 156414 80036
rect 156478 79971 156506 80036
rect 156464 79962 156520 79971
rect 155730 79834 155782 79840
rect 155914 79892 155966 79898
rect 155914 79834 155966 79840
rect 156006 79892 156058 79898
rect 156006 79834 156058 79840
rect 156374 79892 156426 79898
rect 156464 79897 156520 79906
rect 156570 79898 156598 80036
rect 156374 79834 156426 79840
rect 156558 79892 156610 79898
rect 156558 79834 156610 79840
rect 156662 79801 156690 80036
rect 156754 79937 156782 80036
rect 156846 79966 156874 80036
rect 156834 79960 156886 79966
rect 156740 79928 156796 79937
rect 156834 79902 156886 79908
rect 156740 79863 156796 79872
rect 156788 79824 156840 79830
rect 155314 79727 155370 79736
rect 155408 79756 155460 79762
rect 155224 79552 155276 79558
rect 155224 79494 155276 79500
rect 155236 78826 155264 79494
rect 155328 78946 155356 79727
rect 155408 79698 155460 79704
rect 155512 79750 155678 79778
rect 156648 79792 156704 79801
rect 155868 79756 155920 79762
rect 155316 78940 155368 78946
rect 155316 78882 155368 78888
rect 155236 78798 155356 78826
rect 155224 78736 155276 78742
rect 155224 78678 155276 78684
rect 155052 71746 155172 71774
rect 155052 71466 155080 71746
rect 155236 71534 155264 78678
rect 155328 75274 155356 78798
rect 155420 77110 155448 79698
rect 155408 77104 155460 77110
rect 155408 77046 155460 77052
rect 155316 75268 155368 75274
rect 155316 75210 155368 75216
rect 155512 74390 155540 79750
rect 155868 79698 155920 79704
rect 156236 79756 156288 79762
rect 156788 79766 156840 79772
rect 156648 79727 156704 79736
rect 156236 79698 156288 79704
rect 155684 79688 155736 79694
rect 155684 79630 155736 79636
rect 155696 75721 155724 79630
rect 155776 79552 155828 79558
rect 155776 79494 155828 79500
rect 155682 75712 155738 75721
rect 155682 75647 155738 75656
rect 155500 74384 155552 74390
rect 155500 74326 155552 74332
rect 155224 71528 155276 71534
rect 155224 71470 155276 71476
rect 155040 71460 155092 71466
rect 155040 71402 155092 71408
rect 154684 70366 154988 70394
rect 154684 69494 154712 70366
rect 155788 69970 155816 79494
rect 155880 73914 155908 79698
rect 156144 79620 156196 79626
rect 156144 79562 156196 79568
rect 156156 77518 156184 79562
rect 156144 77512 156196 77518
rect 156144 77454 156196 77460
rect 155868 73908 155920 73914
rect 155868 73850 155920 73856
rect 156248 73710 156276 79698
rect 156328 79620 156380 79626
rect 156328 79562 156380 79568
rect 156512 79620 156564 79626
rect 156512 79562 156564 79568
rect 156236 73704 156288 73710
rect 156236 73646 156288 73652
rect 156340 73098 156368 79562
rect 156420 79552 156472 79558
rect 156420 79494 156472 79500
rect 156432 76430 156460 79494
rect 156420 76424 156472 76430
rect 156420 76366 156472 76372
rect 156328 73092 156380 73098
rect 156328 73034 156380 73040
rect 155960 72480 156012 72486
rect 155960 72422 156012 72428
rect 155776 69964 155828 69970
rect 155776 69906 155828 69912
rect 154672 69488 154724 69494
rect 154672 69430 154724 69436
rect 154040 64846 154252 64874
rect 154040 28966 154068 64846
rect 154028 28960 154080 28966
rect 154028 28902 154080 28908
rect 153936 23044 153988 23050
rect 153936 22986 153988 22992
rect 153844 22976 153896 22982
rect 153844 22918 153896 22924
rect 153660 20324 153712 20330
rect 153660 20266 153712 20272
rect 155972 16574 156000 72422
rect 156524 70394 156552 79562
rect 156604 79552 156656 79558
rect 156604 79494 156656 79500
rect 156616 71398 156644 79494
rect 156694 78976 156750 78985
rect 156694 78911 156750 78920
rect 156708 76498 156736 78911
rect 156696 76492 156748 76498
rect 156696 76434 156748 76440
rect 156800 75585 156828 79766
rect 156938 79336 156966 80036
rect 157030 79801 157058 80036
rect 157122 79966 157150 80036
rect 157214 79966 157242 80036
rect 157110 79960 157162 79966
rect 157110 79902 157162 79908
rect 157202 79960 157254 79966
rect 157202 79902 157254 79908
rect 157306 79898 157334 80036
rect 157398 79966 157426 80036
rect 157490 79966 157518 80036
rect 157582 79966 157610 80036
rect 157674 79966 157702 80036
rect 157766 79971 157794 80036
rect 157386 79960 157438 79966
rect 157386 79902 157438 79908
rect 157478 79960 157530 79966
rect 157478 79902 157530 79908
rect 157570 79960 157622 79966
rect 157570 79902 157622 79908
rect 157662 79960 157714 79966
rect 157662 79902 157714 79908
rect 157752 79962 157808 79971
rect 157294 79892 157346 79898
rect 157752 79897 157808 79906
rect 157858 79898 157886 80036
rect 157950 79971 157978 80036
rect 157936 79962 157992 79971
rect 157294 79834 157346 79840
rect 157846 79892 157898 79898
rect 157936 79897 157992 79906
rect 158042 79898 158070 80036
rect 157846 79834 157898 79840
rect 158030 79892 158082 79898
rect 158030 79834 158082 79840
rect 158134 79830 158162 80036
rect 158226 79898 158254 80036
rect 158318 79966 158346 80036
rect 158410 79966 158438 80036
rect 158306 79960 158358 79966
rect 158306 79902 158358 79908
rect 158398 79960 158450 79966
rect 158502 79937 158530 80036
rect 158594 79966 158622 80036
rect 158686 79966 158714 80036
rect 158582 79960 158634 79966
rect 158398 79902 158450 79908
rect 158488 79928 158544 79937
rect 158214 79892 158266 79898
rect 158582 79902 158634 79908
rect 158674 79960 158726 79966
rect 158674 79902 158726 79908
rect 158488 79863 158544 79872
rect 158214 79834 158266 79840
rect 158122 79824 158174 79830
rect 157016 79792 157072 79801
rect 158122 79766 158174 79772
rect 158352 79824 158404 79830
rect 158352 79766 158404 79772
rect 158444 79824 158496 79830
rect 158582 79824 158634 79830
rect 158444 79766 158496 79772
rect 158580 79792 158582 79801
rect 158634 79792 158636 79801
rect 157016 79727 157072 79736
rect 157156 79756 157208 79762
rect 157156 79698 157208 79704
rect 158260 79756 158312 79762
rect 158260 79698 158312 79704
rect 157064 79552 157116 79558
rect 157064 79494 157116 79500
rect 157076 79370 157104 79494
rect 156892 79308 156966 79336
rect 157030 79342 157104 79370
rect 156786 75576 156842 75585
rect 156786 75511 156842 75520
rect 156892 75449 156920 79308
rect 157030 79200 157058 79342
rect 157030 79172 157104 79200
rect 156970 75984 157026 75993
rect 156970 75919 157026 75928
rect 156878 75440 156934 75449
rect 156878 75375 156934 75384
rect 156880 75268 156932 75274
rect 156880 75210 156932 75216
rect 156604 71392 156656 71398
rect 156604 71334 156656 71340
rect 156064 70366 156552 70394
rect 156064 70310 156092 70366
rect 156052 70304 156104 70310
rect 156052 70246 156104 70252
rect 156892 68814 156920 75210
rect 156984 70106 157012 75919
rect 157076 74050 157104 79172
rect 157168 76129 157196 79698
rect 157248 79688 157300 79694
rect 157248 79630 157300 79636
rect 157616 79688 157668 79694
rect 158168 79688 158220 79694
rect 157616 79630 157668 79636
rect 157706 79656 157762 79665
rect 157154 76120 157210 76129
rect 157154 76055 157210 76064
rect 157064 74044 157116 74050
rect 157064 73986 157116 73992
rect 157260 73953 157288 79630
rect 157340 79620 157392 79626
rect 157340 79562 157392 79568
rect 157524 79620 157576 79626
rect 157524 79562 157576 79568
rect 157352 78742 157380 79562
rect 157432 79212 157484 79218
rect 157432 79154 157484 79160
rect 157444 79121 157472 79154
rect 157430 79112 157486 79121
rect 157430 79047 157486 79056
rect 157340 78736 157392 78742
rect 157340 78678 157392 78684
rect 157536 76158 157564 79562
rect 157524 76152 157576 76158
rect 157524 76094 157576 76100
rect 157628 74458 157656 79630
rect 158168 79630 158220 79636
rect 157706 79591 157762 79600
rect 157800 79620 157852 79626
rect 157720 75614 157748 79591
rect 157800 79562 157852 79568
rect 157812 78198 157840 79562
rect 157984 79552 158036 79558
rect 157904 79512 157984 79540
rect 157800 78192 157852 78198
rect 157800 78134 157852 78140
rect 157904 77450 157932 79512
rect 157984 79494 158036 79500
rect 158076 79416 158128 79422
rect 158076 79358 158128 79364
rect 158088 79150 158116 79358
rect 158076 79144 158128 79150
rect 158076 79086 158128 79092
rect 157892 77444 157944 77450
rect 157892 77386 157944 77392
rect 157708 75608 157760 75614
rect 157708 75550 157760 75556
rect 157708 75336 157760 75342
rect 157708 75278 157760 75284
rect 157616 74452 157668 74458
rect 157616 74394 157668 74400
rect 157614 74352 157670 74361
rect 157614 74287 157670 74296
rect 157628 74254 157656 74287
rect 157616 74248 157668 74254
rect 157616 74190 157668 74196
rect 157246 73944 157302 73953
rect 157246 73879 157302 73888
rect 157614 73808 157670 73817
rect 157614 73743 157616 73752
rect 157668 73743 157670 73752
rect 157616 73714 157668 73720
rect 156972 70100 157024 70106
rect 156972 70042 157024 70048
rect 157720 70038 157748 75278
rect 158180 73642 158208 79630
rect 158272 76378 158300 79698
rect 158364 79665 158392 79766
rect 158350 79656 158406 79665
rect 158350 79591 158406 79600
rect 158352 79484 158404 79490
rect 158352 79426 158404 79432
rect 158364 79014 158392 79426
rect 158352 79008 158404 79014
rect 158352 78950 158404 78956
rect 158456 77058 158484 79766
rect 158778 79778 158806 80036
rect 158870 79898 158898 80036
rect 158962 79898 158990 80036
rect 158858 79892 158910 79898
rect 158858 79834 158910 79840
rect 158950 79892 159002 79898
rect 158950 79834 159002 79840
rect 159054 79812 159082 80036
rect 159146 79966 159174 80036
rect 159238 79966 159266 80036
rect 159134 79960 159186 79966
rect 159134 79902 159186 79908
rect 159226 79960 159278 79966
rect 159330 79937 159358 80036
rect 159226 79902 159278 79908
rect 159316 79928 159372 79937
rect 159316 79863 159372 79872
rect 159054 79784 159312 79812
rect 158778 79750 158852 79778
rect 158580 79727 158636 79736
rect 158628 79688 158680 79694
rect 158680 79648 158760 79676
rect 158628 79630 158680 79636
rect 158628 79484 158680 79490
rect 158628 79426 158680 79432
rect 158536 79416 158588 79422
rect 158536 79358 158588 79364
rect 158548 78810 158576 79358
rect 158640 78985 158668 79426
rect 158626 78976 158682 78985
rect 158626 78911 158682 78920
rect 158536 78804 158588 78810
rect 158536 78746 158588 78752
rect 158732 78402 158760 79648
rect 158824 78878 158852 79750
rect 159180 79688 159232 79694
rect 159284 79665 159312 79784
rect 159422 79744 159450 80036
rect 159514 79966 159542 80036
rect 159502 79960 159554 79966
rect 159502 79902 159554 79908
rect 159606 79744 159634 80036
rect 159698 79966 159726 80036
rect 159790 79966 159818 80036
rect 159686 79960 159738 79966
rect 159686 79902 159738 79908
rect 159778 79960 159830 79966
rect 159778 79902 159830 79908
rect 159882 79744 159910 80036
rect 159974 79812 160002 80036
rect 160066 79966 160094 80036
rect 160158 79966 160186 80036
rect 160250 79966 160278 80036
rect 160054 79960 160106 79966
rect 160054 79902 160106 79908
rect 160146 79960 160198 79966
rect 160146 79902 160198 79908
rect 160238 79960 160290 79966
rect 160238 79902 160290 79908
rect 160342 79898 160370 80036
rect 160434 79966 160462 80036
rect 160526 79971 160554 80036
rect 160422 79960 160474 79966
rect 160422 79902 160474 79908
rect 160512 79962 160568 79971
rect 160618 79966 160646 80036
rect 160330 79892 160382 79898
rect 160512 79897 160568 79906
rect 160606 79960 160658 79966
rect 160606 79902 160658 79908
rect 160330 79834 160382 79840
rect 160468 79824 160520 79830
rect 159974 79784 160048 79812
rect 159422 79716 159496 79744
rect 159606 79716 159772 79744
rect 159882 79716 159956 79744
rect 159180 79630 159232 79636
rect 159270 79656 159326 79665
rect 158996 79620 159048 79626
rect 158996 79562 159048 79568
rect 159088 79620 159140 79626
rect 159088 79562 159140 79568
rect 158904 79552 158956 79558
rect 158904 79494 158956 79500
rect 158812 78872 158864 78878
rect 158812 78814 158864 78820
rect 158720 78396 158772 78402
rect 158720 78338 158772 78344
rect 158812 77444 158864 77450
rect 158812 77386 158864 77392
rect 158456 77030 158668 77058
rect 158442 76936 158498 76945
rect 158442 76871 158498 76880
rect 158272 76350 158392 76378
rect 158258 76256 158314 76265
rect 158258 76191 158314 76200
rect 158168 73636 158220 73642
rect 158168 73578 158220 73584
rect 157708 70032 157760 70038
rect 157708 69974 157760 69980
rect 156880 68808 156932 68814
rect 156880 68750 156932 68756
rect 158272 67046 158300 76191
rect 158364 72690 158392 76350
rect 158456 73982 158484 76871
rect 158536 75948 158588 75954
rect 158536 75890 158588 75896
rect 158444 73976 158496 73982
rect 158444 73918 158496 73924
rect 158352 72684 158404 72690
rect 158352 72626 158404 72632
rect 158548 70174 158576 75890
rect 158640 73817 158668 77030
rect 158824 74534 158852 77386
rect 158916 76702 158944 79494
rect 158904 76696 158956 76702
rect 158904 76638 158956 76644
rect 158824 74506 158944 74534
rect 158626 73808 158682 73817
rect 158626 73743 158682 73752
rect 158916 71330 158944 74506
rect 159008 72758 159036 79562
rect 158996 72752 159048 72758
rect 158996 72694 159048 72700
rect 159100 72282 159128 79562
rect 159192 75410 159220 79630
rect 159270 79591 159326 79600
rect 159272 79552 159324 79558
rect 159272 79494 159324 79500
rect 159180 75404 159232 75410
rect 159180 75346 159232 75352
rect 159284 72554 159312 79494
rect 159364 79212 159416 79218
rect 159364 79154 159416 79160
rect 159376 76974 159404 79154
rect 159364 76968 159416 76974
rect 159364 76910 159416 76916
rect 159468 72826 159496 79716
rect 159638 79656 159694 79665
rect 159548 79620 159600 79626
rect 159638 79591 159694 79600
rect 159548 79562 159600 79568
rect 159560 72894 159588 79562
rect 159548 72888 159600 72894
rect 159548 72830 159600 72836
rect 159456 72820 159508 72826
rect 159456 72762 159508 72768
rect 159272 72548 159324 72554
rect 159272 72490 159324 72496
rect 159088 72276 159140 72282
rect 159088 72218 159140 72224
rect 158904 71324 158956 71330
rect 158904 71266 158956 71272
rect 158536 70168 158588 70174
rect 158536 70110 158588 70116
rect 159652 68678 159680 79591
rect 159744 75954 159772 79716
rect 159824 79620 159876 79626
rect 159824 79562 159876 79568
rect 159732 75948 159784 75954
rect 159732 75890 159784 75896
rect 159836 75614 159864 79562
rect 159928 78130 159956 79716
rect 159916 78124 159968 78130
rect 159916 78066 159968 78072
rect 159916 75948 159968 75954
rect 159916 75890 159968 75896
rect 159732 75608 159784 75614
rect 159732 75550 159784 75556
rect 159824 75608 159876 75614
rect 159824 75550 159876 75556
rect 159744 72962 159772 75550
rect 159732 72956 159784 72962
rect 159732 72898 159784 72904
rect 159928 71194 159956 75890
rect 160020 74905 160048 79784
rect 160710 79812 160738 80036
rect 160802 79966 160830 80036
rect 160894 79966 160922 80036
rect 160790 79960 160842 79966
rect 160790 79902 160842 79908
rect 160882 79960 160934 79966
rect 160986 79937 161014 80036
rect 160882 79902 160934 79908
rect 160972 79928 161028 79937
rect 161078 79898 161106 80036
rect 161170 79898 161198 80036
rect 161262 79966 161290 80036
rect 161354 79971 161382 80036
rect 161250 79960 161302 79966
rect 161250 79902 161302 79908
rect 161340 79962 161396 79971
rect 161446 79966 161474 80036
rect 160972 79863 161028 79872
rect 161066 79892 161118 79898
rect 161066 79834 161118 79840
rect 161158 79892 161210 79898
rect 161340 79897 161396 79906
rect 161434 79960 161486 79966
rect 161434 79902 161486 79908
rect 161158 79834 161210 79840
rect 160468 79766 160520 79772
rect 160664 79784 160738 79812
rect 161110 79792 161166 79801
rect 160192 79688 160244 79694
rect 160480 79642 160508 79766
rect 160560 79756 160612 79762
rect 160560 79698 160612 79704
rect 160192 79630 160244 79636
rect 160100 79212 160152 79218
rect 160100 79154 160152 79160
rect 160112 79014 160140 79154
rect 160100 79008 160152 79014
rect 160100 78950 160152 78956
rect 160098 76936 160154 76945
rect 160098 76871 160154 76880
rect 160006 74896 160062 74905
rect 160006 74831 160062 74840
rect 159916 71188 159968 71194
rect 159916 71130 159968 71136
rect 159640 68672 159692 68678
rect 159640 68614 159692 68620
rect 158260 67040 158312 67046
rect 158260 66982 158312 66988
rect 155972 16546 156184 16574
rect 153568 14952 153620 14958
rect 153568 14894 153620 14900
rect 153476 6520 153528 6526
rect 153476 6462 153528 6468
rect 153384 6452 153436 6458
rect 153384 6394 153436 6400
rect 153292 6384 153344 6390
rect 153292 6326 153344 6332
rect 153200 6316 153252 6322
rect 153200 6258 153252 6264
rect 155408 5228 155460 5234
rect 155408 5170 155460 5176
rect 153016 4140 153068 4146
rect 153016 4082 153068 4088
rect 151820 3800 151872 3806
rect 151820 3742 151872 3748
rect 150530 3632 150586 3641
rect 149244 3596 149296 3602
rect 150530 3567 150586 3576
rect 149244 3538 149296 3544
rect 149072 3454 149560 3482
rect 149532 480 149560 3454
rect 150624 3188 150676 3194
rect 150624 3130 150676 3136
rect 150636 480 150664 3130
rect 151832 480 151860 3742
rect 153028 480 153056 4082
rect 154212 3052 154264 3058
rect 154212 2994 154264 3000
rect 154224 480 154252 2994
rect 155420 480 155448 5170
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 160112 14890 160140 76871
rect 160204 75070 160232 79630
rect 160388 79614 160508 79642
rect 160284 79552 160336 79558
rect 160284 79494 160336 79500
rect 160296 76838 160324 79494
rect 160388 77450 160416 79614
rect 160468 79552 160520 79558
rect 160468 79494 160520 79500
rect 160376 77444 160428 77450
rect 160376 77386 160428 77392
rect 160284 76832 160336 76838
rect 160284 76774 160336 76780
rect 160284 76628 160336 76634
rect 160284 76570 160336 76576
rect 160192 75064 160244 75070
rect 160192 75006 160244 75012
rect 160296 74882 160324 76570
rect 160376 76084 160428 76090
rect 160376 76026 160428 76032
rect 160204 74854 160324 74882
rect 160100 14884 160152 14890
rect 160100 14826 160152 14832
rect 160204 14822 160232 74854
rect 160284 74792 160336 74798
rect 160284 74734 160336 74740
rect 160192 14816 160244 14822
rect 160192 14758 160244 14764
rect 160296 14754 160324 74734
rect 160388 26926 160416 76026
rect 160480 31618 160508 79494
rect 160572 76090 160600 79698
rect 160664 76770 160692 79784
rect 161110 79727 161166 79736
rect 161296 79756 161348 79762
rect 160744 79688 160796 79694
rect 161124 79676 161152 79727
rect 161538 79744 161566 80036
rect 161630 79937 161658 80036
rect 161722 79966 161750 80036
rect 161710 79960 161762 79966
rect 161616 79928 161672 79937
rect 161710 79902 161762 79908
rect 161616 79863 161672 79872
rect 161814 79830 161842 80036
rect 161906 79898 161934 80036
rect 161998 79971 162026 80036
rect 161984 79962 162040 79971
rect 162090 79966 162118 80036
rect 161894 79892 161946 79898
rect 161984 79897 162040 79906
rect 162078 79960 162130 79966
rect 162078 79902 162130 79908
rect 161894 79834 161946 79840
rect 161802 79824 161854 79830
rect 162182 79812 162210 80036
rect 162274 79830 162302 80036
rect 162366 79971 162394 80036
rect 162352 79962 162408 79971
rect 162352 79897 162408 79906
rect 161802 79766 161854 79772
rect 162136 79784 162210 79812
rect 162262 79824 162314 79830
rect 161296 79698 161348 79704
rect 161492 79716 161566 79744
rect 161664 79756 161716 79762
rect 160744 79630 160796 79636
rect 161032 79648 161152 79676
rect 161202 79656 161258 79665
rect 160652 76764 160704 76770
rect 160652 76706 160704 76712
rect 160756 76634 160784 79630
rect 160836 79620 160888 79626
rect 160836 79562 160888 79568
rect 160744 76628 160796 76634
rect 160744 76570 160796 76576
rect 160560 76084 160612 76090
rect 160560 76026 160612 76032
rect 160848 75970 160876 79562
rect 160928 79552 160980 79558
rect 160928 79494 160980 79500
rect 160572 75942 160876 75970
rect 160468 31612 160520 31618
rect 160468 31554 160520 31560
rect 160572 31550 160600 75942
rect 160652 75064 160704 75070
rect 160652 75006 160704 75012
rect 160664 64258 160692 75006
rect 160940 74798 160968 79494
rect 161032 78674 161060 79648
rect 161202 79591 161258 79600
rect 161112 79552 161164 79558
rect 161112 79494 161164 79500
rect 161124 78849 161152 79494
rect 161110 78840 161166 78849
rect 161110 78775 161166 78784
rect 161216 78742 161244 79591
rect 161112 78736 161164 78742
rect 161112 78678 161164 78684
rect 161204 78736 161256 78742
rect 161204 78678 161256 78684
rect 161020 78668 161072 78674
rect 161020 78610 161072 78616
rect 160928 74792 160980 74798
rect 160928 74734 160980 74740
rect 161124 74118 161152 78678
rect 161308 77353 161336 79698
rect 161492 79608 161520 79716
rect 161664 79698 161716 79704
rect 161400 79580 161520 79608
rect 161400 78334 161428 79580
rect 161572 79552 161624 79558
rect 161572 79494 161624 79500
rect 161480 79484 161532 79490
rect 161480 79426 161532 79432
rect 161388 78328 161440 78334
rect 161388 78270 161440 78276
rect 161294 77344 161350 77353
rect 161294 77279 161350 77288
rect 161112 74112 161164 74118
rect 161112 74054 161164 74060
rect 160652 64252 160704 64258
rect 160652 64194 160704 64200
rect 160560 31544 160612 31550
rect 160560 31486 160612 31492
rect 160376 26920 160428 26926
rect 160376 26862 160428 26868
rect 160284 14748 160336 14754
rect 160284 14690 160336 14696
rect 161492 9042 161520 79426
rect 161584 78849 161612 79494
rect 161570 78840 161626 78849
rect 161676 78826 161704 79698
rect 162032 79552 162084 79558
rect 162032 79494 162084 79500
rect 161938 78840 161994 78849
rect 161676 78798 161796 78826
rect 161570 78775 161626 78784
rect 161572 78464 161624 78470
rect 161572 78406 161624 78412
rect 161584 75154 161612 78406
rect 161664 78260 161716 78266
rect 161664 78202 161716 78208
rect 161676 75274 161704 78202
rect 161664 75268 161716 75274
rect 161664 75210 161716 75216
rect 161584 75126 161704 75154
rect 161572 75064 161624 75070
rect 161572 75006 161624 75012
rect 161584 11898 161612 75006
rect 161676 11966 161704 75126
rect 161768 14686 161796 78798
rect 161938 78775 161994 78784
rect 161846 78704 161902 78713
rect 161846 78639 161902 78648
rect 161860 76566 161888 78639
rect 161848 76560 161900 76566
rect 161848 76502 161900 76508
rect 161848 75268 161900 75274
rect 161848 75210 161900 75216
rect 161860 17610 161888 75210
rect 161952 20262 161980 78775
rect 162044 78470 162072 79494
rect 162032 78464 162084 78470
rect 162032 78406 162084 78412
rect 162136 75070 162164 79784
rect 162458 79801 162486 80036
rect 162550 79966 162578 80036
rect 162538 79960 162590 79966
rect 162538 79902 162590 79908
rect 162262 79766 162314 79772
rect 162444 79792 162500 79801
rect 162444 79727 162500 79736
rect 162400 79688 162452 79694
rect 162400 79630 162452 79636
rect 162216 79620 162268 79626
rect 162216 79562 162268 79568
rect 162228 77926 162256 79562
rect 162306 78976 162362 78985
rect 162306 78911 162362 78920
rect 162216 77920 162268 77926
rect 162216 77862 162268 77868
rect 162124 75064 162176 75070
rect 162124 75006 162176 75012
rect 162320 70394 162348 78911
rect 162412 78810 162440 79630
rect 162642 79608 162670 80036
rect 162734 79971 162762 80036
rect 162720 79962 162776 79971
rect 162826 79966 162854 80036
rect 162918 79966 162946 80036
rect 162720 79897 162776 79906
rect 162814 79960 162866 79966
rect 162814 79902 162866 79908
rect 162906 79960 162958 79966
rect 162906 79902 162958 79908
rect 163010 79830 163038 80036
rect 162814 79824 162866 79830
rect 162814 79766 162866 79772
rect 162998 79824 163050 79830
rect 162998 79766 163050 79772
rect 162826 79676 162854 79766
rect 163102 79744 163130 80036
rect 163194 79937 163222 80036
rect 163180 79928 163236 79937
rect 163180 79863 163236 79872
rect 163286 79744 163314 80036
rect 163102 79716 163176 79744
rect 162826 79648 162946 79676
rect 162596 79580 162670 79608
rect 162492 79484 162544 79490
rect 162492 79426 162544 79432
rect 162400 78804 162452 78810
rect 162400 78746 162452 78752
rect 162504 78713 162532 79426
rect 162596 79014 162624 79580
rect 162918 79540 162946 79648
rect 162872 79512 162946 79540
rect 162768 79484 162820 79490
rect 162768 79426 162820 79432
rect 162584 79008 162636 79014
rect 162584 78950 162636 78956
rect 162584 78736 162636 78742
rect 162490 78704 162546 78713
rect 162400 78668 162452 78674
rect 162584 78678 162636 78684
rect 162676 78736 162728 78742
rect 162676 78678 162728 78684
rect 162490 78639 162546 78648
rect 162400 78610 162452 78616
rect 162136 70366 162348 70394
rect 162412 70394 162440 78610
rect 162412 70366 162532 70394
rect 162136 64874 162164 70366
rect 162044 64846 162164 64874
rect 162044 28762 162072 64846
rect 162032 28756 162084 28762
rect 162032 28698 162084 28704
rect 162504 25906 162532 70366
rect 162596 25974 162624 78678
rect 162688 78266 162716 78678
rect 162676 78260 162728 78266
rect 162676 78202 162728 78208
rect 162780 77294 162808 79426
rect 162872 79121 162900 79512
rect 163044 79484 163096 79490
rect 163044 79426 163096 79432
rect 162858 79112 162914 79121
rect 162858 79047 162914 79056
rect 162860 79008 162912 79014
rect 162860 78950 162912 78956
rect 162872 77994 162900 78950
rect 162860 77988 162912 77994
rect 162860 77930 162912 77936
rect 162780 77266 162992 77294
rect 162860 75200 162912 75206
rect 162860 75142 162912 75148
rect 162584 25968 162636 25974
rect 162584 25910 162636 25916
rect 162492 25900 162544 25906
rect 162492 25842 162544 25848
rect 161940 20256 161992 20262
rect 161940 20198 161992 20204
rect 161848 17604 161900 17610
rect 161848 17546 161900 17552
rect 161756 14680 161808 14686
rect 161756 14622 161808 14628
rect 162872 14618 162900 75142
rect 162964 28694 162992 77266
rect 163056 31482 163084 79426
rect 163148 75274 163176 79716
rect 163240 79716 163314 79744
rect 163378 79744 163406 80036
rect 163470 79898 163498 80036
rect 163562 79898 163590 80036
rect 163654 79971 163682 80036
rect 163640 79962 163696 79971
rect 163458 79892 163510 79898
rect 163458 79834 163510 79840
rect 163550 79892 163602 79898
rect 163640 79897 163696 79906
rect 163746 79898 163774 80036
rect 163838 79966 163866 80036
rect 163930 79966 163958 80036
rect 163826 79960 163878 79966
rect 163826 79902 163878 79908
rect 163918 79960 163970 79966
rect 163918 79902 163970 79908
rect 163550 79834 163602 79840
rect 163734 79892 163786 79898
rect 163734 79834 163786 79840
rect 164022 79830 164050 80036
rect 164114 79937 164142 80036
rect 164100 79928 164156 79937
rect 164100 79863 164156 79872
rect 164010 79824 164062 79830
rect 164206 79812 164234 80036
rect 164298 79898 164326 80036
rect 164390 79971 164418 80036
rect 164376 79962 164432 79971
rect 164482 79966 164510 80036
rect 164286 79892 164338 79898
rect 164376 79897 164432 79906
rect 164470 79960 164522 79966
rect 164470 79902 164522 79908
rect 164574 79898 164602 80036
rect 164286 79834 164338 79840
rect 164562 79892 164614 79898
rect 164562 79834 164614 79840
rect 164010 79766 164062 79772
rect 164160 79784 164234 79812
rect 163504 79756 163556 79762
rect 163378 79716 163452 79744
rect 163240 79014 163268 79716
rect 163228 79008 163280 79014
rect 163228 78950 163280 78956
rect 163424 78826 163452 79716
rect 163504 79698 163556 79704
rect 163516 79490 163544 79698
rect 163596 79688 163648 79694
rect 163594 79656 163596 79665
rect 163688 79688 163740 79694
rect 163648 79656 163650 79665
rect 163688 79630 163740 79636
rect 163964 79688 164016 79694
rect 163964 79630 164016 79636
rect 163594 79591 163650 79600
rect 163504 79484 163556 79490
rect 163504 79426 163556 79432
rect 163502 79112 163558 79121
rect 163502 79047 163558 79056
rect 163240 78798 163452 78826
rect 163136 75268 163188 75274
rect 163136 75210 163188 75216
rect 163240 75206 163268 78798
rect 163318 78704 163374 78713
rect 163318 78639 163374 78648
rect 163228 75200 163280 75206
rect 163228 75142 163280 75148
rect 163136 75132 163188 75138
rect 163136 75074 163188 75080
rect 163044 31476 163096 31482
rect 163044 31418 163096 31424
rect 163148 31414 163176 75074
rect 163228 75064 163280 75070
rect 163228 75006 163280 75012
rect 163240 34134 163268 75006
rect 163332 34270 163360 78639
rect 163516 77294 163544 79047
rect 163596 79008 163648 79014
rect 163596 78950 163648 78956
rect 163424 77266 163544 77294
rect 163320 34264 163372 34270
rect 163320 34206 163372 34212
rect 163424 34202 163452 77266
rect 163608 76945 163636 78950
rect 163700 77314 163728 79630
rect 163780 79620 163832 79626
rect 163780 79562 163832 79568
rect 163872 79620 163924 79626
rect 163872 79562 163924 79568
rect 163688 77308 163740 77314
rect 163688 77250 163740 77256
rect 163594 76936 163650 76945
rect 163594 76871 163650 76880
rect 163504 75268 163556 75274
rect 163504 75210 163556 75216
rect 163516 34338 163544 75210
rect 163792 75138 163820 79562
rect 163780 75132 163832 75138
rect 163780 75074 163832 75080
rect 163884 75070 163912 79562
rect 163976 78713 164004 79630
rect 164056 79620 164108 79626
rect 164056 79562 164108 79568
rect 164068 79150 164096 79562
rect 164056 79144 164108 79150
rect 164056 79086 164108 79092
rect 164054 78976 164110 78985
rect 164054 78911 164110 78920
rect 163962 78704 164018 78713
rect 163962 78639 164018 78648
rect 164068 78470 164096 78911
rect 164160 78849 164188 79784
rect 164332 79756 164384 79762
rect 164332 79698 164384 79704
rect 164240 79620 164292 79626
rect 164240 79562 164292 79568
rect 164146 78840 164202 78849
rect 164146 78775 164202 78784
rect 164252 78674 164280 79562
rect 164240 78668 164292 78674
rect 164240 78610 164292 78616
rect 164056 78464 164108 78470
rect 164056 78406 164108 78412
rect 163964 78396 164016 78402
rect 163964 78338 164016 78344
rect 163872 75064 163924 75070
rect 163872 75006 163924 75012
rect 163976 64874 164004 78338
rect 164344 77382 164372 79698
rect 164666 79676 164694 80036
rect 164758 79937 164786 80036
rect 164744 79928 164800 79937
rect 164744 79863 164800 79872
rect 164850 79744 164878 80036
rect 164942 79898 164970 80036
rect 165034 79898 165062 80036
rect 165126 79898 165154 80036
rect 165218 79937 165246 80036
rect 165204 79928 165260 79937
rect 164930 79892 164982 79898
rect 164930 79834 164982 79840
rect 165022 79892 165074 79898
rect 165022 79834 165074 79840
rect 165114 79892 165166 79898
rect 165310 79898 165338 80036
rect 165204 79863 165260 79872
rect 165298 79892 165350 79898
rect 165114 79834 165166 79840
rect 165298 79834 165350 79840
rect 164514 79656 164570 79665
rect 164514 79591 164570 79600
rect 164620 79648 164694 79676
rect 164804 79716 164878 79744
rect 164976 79756 165028 79762
rect 164424 79552 164476 79558
rect 164424 79494 164476 79500
rect 164436 78985 164464 79494
rect 164528 79082 164556 79591
rect 164516 79076 164568 79082
rect 164516 79018 164568 79024
rect 164422 78976 164478 78985
rect 164422 78911 164478 78920
rect 164620 78674 164648 79648
rect 164700 79552 164752 79558
rect 164700 79494 164752 79500
rect 164424 78668 164476 78674
rect 164424 78610 164476 78616
rect 164608 78668 164660 78674
rect 164608 78610 164660 78616
rect 164332 77376 164384 77382
rect 164332 77318 164384 77324
rect 164332 75336 164384 75342
rect 164332 75278 164384 75284
rect 164240 75132 164292 75138
rect 164240 75074 164292 75080
rect 163884 64846 164004 64874
rect 163884 34406 163912 64846
rect 163872 34400 163924 34406
rect 163872 34342 163924 34348
rect 163504 34332 163556 34338
rect 163504 34274 163556 34280
rect 163412 34196 163464 34202
rect 163412 34138 163464 34144
rect 163228 34128 163280 34134
rect 163228 34070 163280 34076
rect 163136 31408 163188 31414
rect 163136 31350 163188 31356
rect 162952 28688 163004 28694
rect 162952 28630 163004 28636
rect 162950 18728 163006 18737
rect 162950 18663 163006 18672
rect 162964 16574 162992 18663
rect 162964 16546 163728 16574
rect 162860 14612 162912 14618
rect 162860 14554 162912 14560
rect 161664 11960 161716 11966
rect 161664 11902 161716 11908
rect 161572 11892 161624 11898
rect 161572 11834 161624 11840
rect 161480 9036 161532 9042
rect 161480 8978 161532 8984
rect 157800 5160 157852 5166
rect 157800 5102 157852 5108
rect 156696 4072 156748 4078
rect 156696 4014 156748 4020
rect 156708 3398 156736 4014
rect 156696 3392 156748 3398
rect 156696 3334 156748 3340
rect 157812 480 157840 5102
rect 162490 4992 162546 5001
rect 162490 4927 162546 4936
rect 158904 4888 158956 4894
rect 158904 4830 158956 4836
rect 158916 480 158944 4830
rect 160100 3868 160152 3874
rect 160100 3810 160152 3816
rect 160112 480 160140 3810
rect 161296 3732 161348 3738
rect 161296 3674 161348 3680
rect 161308 480 161336 3674
rect 162504 480 162532 4927
rect 163700 480 163728 16546
rect 164252 7614 164280 75074
rect 164344 17474 164372 75278
rect 164436 17542 164464 78610
rect 164608 78192 164660 78198
rect 164608 78134 164660 78140
rect 164620 76362 164648 78134
rect 164608 76356 164660 76362
rect 164608 76298 164660 76304
rect 164516 75268 164568 75274
rect 164516 75210 164568 75216
rect 164528 31346 164556 75210
rect 164608 75200 164660 75206
rect 164608 75142 164660 75148
rect 164620 58750 164648 75142
rect 164712 65550 164740 79494
rect 164804 78810 164832 79716
rect 164976 79698 165028 79704
rect 165160 79756 165212 79762
rect 165160 79698 165212 79704
rect 165252 79756 165304 79762
rect 165402 79744 165430 80036
rect 165494 79937 165522 80036
rect 165480 79928 165536 79937
rect 165480 79863 165536 79872
rect 165586 79830 165614 80036
rect 165678 79898 165706 80036
rect 165770 79966 165798 80036
rect 165758 79960 165810 79966
rect 165758 79902 165810 79908
rect 165666 79892 165718 79898
rect 165666 79834 165718 79840
rect 165574 79824 165626 79830
rect 165862 79812 165890 80036
rect 165954 79966 165982 80036
rect 166046 79966 166074 80036
rect 166138 79966 166166 80036
rect 165942 79960 165994 79966
rect 165942 79902 165994 79908
rect 166034 79960 166086 79966
rect 166034 79902 166086 79908
rect 166126 79960 166178 79966
rect 166126 79902 166178 79908
rect 166230 79830 166258 80036
rect 165988 79824 166040 79830
rect 165862 79784 165936 79812
rect 165574 79766 165626 79772
rect 165712 79756 165764 79762
rect 165402 79716 165476 79744
rect 165252 79698 165304 79704
rect 164884 79076 164936 79082
rect 164884 79018 164936 79024
rect 164792 78804 164844 78810
rect 164792 78746 164844 78752
rect 164792 78668 164844 78674
rect 164792 78610 164844 78616
rect 164804 66910 164832 78610
rect 164896 75274 164924 79018
rect 164884 75268 164936 75274
rect 164884 75210 164936 75216
rect 164988 75206 165016 79698
rect 165068 79688 165120 79694
rect 165068 79630 165120 79636
rect 165080 75342 165108 79630
rect 165068 75336 165120 75342
rect 165068 75278 165120 75284
rect 164976 75200 165028 75206
rect 164976 75142 165028 75148
rect 165172 75138 165200 79698
rect 165264 78713 165292 79698
rect 165250 78704 165306 78713
rect 165250 78639 165306 78648
rect 165448 78033 165476 79716
rect 165712 79698 165764 79704
rect 165528 79688 165580 79694
rect 165528 79630 165580 79636
rect 165540 78713 165568 79630
rect 165620 79416 165672 79422
rect 165620 79358 165672 79364
rect 165632 79121 165660 79358
rect 165618 79112 165674 79121
rect 165618 79047 165674 79056
rect 165526 78704 165582 78713
rect 165724 78656 165752 79698
rect 165804 79688 165856 79694
rect 165804 79630 165856 79636
rect 165816 79218 165844 79630
rect 165908 79506 165936 79784
rect 165988 79766 166040 79772
rect 166080 79824 166132 79830
rect 166080 79766 166132 79772
rect 166218 79824 166270 79830
rect 166218 79766 166270 79772
rect 166000 79626 166028 79766
rect 165988 79620 166040 79626
rect 165988 79562 166040 79568
rect 165908 79478 166028 79506
rect 165896 79416 165948 79422
rect 165896 79358 165948 79364
rect 165804 79212 165856 79218
rect 165804 79154 165856 79160
rect 165526 78639 165582 78648
rect 165632 78628 165752 78656
rect 165434 78024 165490 78033
rect 165434 77959 165490 77968
rect 165436 77444 165488 77450
rect 165436 77386 165488 77392
rect 165344 77308 165396 77314
rect 165344 77250 165396 77256
rect 165252 76356 165304 76362
rect 165252 76298 165304 76304
rect 165160 75132 165212 75138
rect 165160 75074 165212 75080
rect 165160 74996 165212 75002
rect 165160 74938 165212 74944
rect 164792 66904 164844 66910
rect 164792 66846 164844 66852
rect 164700 65544 164752 65550
rect 164700 65486 164752 65492
rect 164608 58744 164660 58750
rect 164608 58686 164660 58692
rect 164516 31340 164568 31346
rect 164516 31282 164568 31288
rect 164424 17536 164476 17542
rect 164424 17478 164476 17484
rect 164332 17468 164384 17474
rect 164332 17410 164384 17416
rect 165172 12034 165200 74938
rect 165264 72622 165292 76298
rect 165252 72616 165304 72622
rect 165252 72558 165304 72564
rect 165356 69834 165384 77250
rect 165448 75002 165476 77386
rect 165632 75274 165660 78628
rect 165908 78520 165936 79358
rect 165724 78492 165936 78520
rect 165620 75268 165672 75274
rect 165620 75210 165672 75216
rect 165436 74996 165488 75002
rect 165436 74938 165488 74944
rect 165344 69828 165396 69834
rect 165344 69770 165396 69776
rect 165160 12028 165212 12034
rect 165160 11970 165212 11976
rect 165724 11830 165752 78492
rect 165804 78124 165856 78130
rect 165804 78066 165856 78072
rect 165816 77314 165844 78066
rect 165804 77308 165856 77314
rect 165804 77250 165856 77256
rect 165896 75336 165948 75342
rect 165896 75278 165948 75284
rect 165804 75200 165856 75206
rect 165804 75142 165856 75148
rect 165816 14550 165844 75142
rect 165908 17406 165936 75278
rect 166000 28558 166028 79478
rect 165988 28552 166040 28558
rect 165988 28494 166040 28500
rect 166092 28490 166120 79766
rect 166172 79688 166224 79694
rect 166172 79630 166224 79636
rect 166184 78674 166212 79630
rect 166322 79608 166350 80036
rect 166414 79898 166442 80036
rect 166402 79892 166454 79898
rect 166402 79834 166454 79840
rect 166506 79744 166534 80036
rect 166598 79937 166626 80036
rect 166584 79928 166640 79937
rect 166584 79863 166640 79872
rect 166690 79744 166718 80036
rect 166782 79898 166810 80036
rect 166874 79966 166902 80036
rect 166862 79960 166914 79966
rect 166862 79902 166914 79908
rect 166966 79898 166994 80036
rect 167058 79937 167086 80036
rect 167150 79966 167178 80036
rect 167138 79960 167190 79966
rect 167044 79928 167100 79937
rect 166770 79892 166822 79898
rect 166770 79834 166822 79840
rect 166954 79892 167006 79898
rect 167138 79902 167190 79908
rect 167242 79898 167270 80036
rect 167044 79863 167100 79872
rect 167230 79892 167282 79898
rect 166954 79834 167006 79840
rect 167230 79834 167282 79840
rect 167334 79778 167362 80036
rect 167426 79898 167454 80036
rect 167518 79937 167546 80036
rect 167610 79966 167638 80036
rect 167702 79971 167730 80036
rect 167598 79960 167650 79966
rect 167504 79928 167560 79937
rect 167414 79892 167466 79898
rect 167598 79902 167650 79908
rect 167688 79962 167744 79971
rect 167794 79966 167822 80036
rect 167886 79966 167914 80036
rect 167978 79966 168006 80036
rect 168070 79966 168098 80036
rect 167688 79897 167744 79906
rect 167782 79960 167834 79966
rect 167782 79902 167834 79908
rect 167874 79960 167926 79966
rect 167874 79902 167926 79908
rect 167966 79960 168018 79966
rect 167966 79902 168018 79908
rect 168058 79960 168110 79966
rect 168058 79902 168110 79908
rect 167504 79863 167560 79872
rect 167414 79834 167466 79840
rect 168162 79812 168190 80036
rect 167092 79756 167144 79762
rect 166506 79716 166580 79744
rect 166690 79716 166764 79744
rect 166276 79580 166350 79608
rect 166172 78668 166224 78674
rect 166172 78610 166224 78616
rect 166172 78328 166224 78334
rect 166172 78270 166224 78276
rect 166184 75410 166212 78270
rect 166172 75404 166224 75410
rect 166172 75346 166224 75352
rect 166172 75268 166224 75274
rect 166172 75210 166224 75216
rect 166184 28626 166212 75210
rect 166276 75206 166304 79580
rect 166356 79484 166408 79490
rect 166356 79426 166408 79432
rect 166264 75200 166316 75206
rect 166264 75142 166316 75148
rect 166368 70394 166396 79426
rect 166552 79150 166580 79716
rect 166630 79656 166686 79665
rect 166630 79591 166686 79600
rect 166644 79558 166672 79591
rect 166632 79552 166684 79558
rect 166632 79494 166684 79500
rect 166632 79416 166684 79422
rect 166632 79358 166684 79364
rect 166540 79144 166592 79150
rect 166540 79086 166592 79092
rect 166446 78840 166502 78849
rect 166446 78775 166502 78784
rect 166460 75342 166488 78775
rect 166644 78656 166672 79358
rect 166736 78849 166764 79716
rect 167092 79698 167144 79704
rect 167184 79756 167236 79762
rect 167184 79698 167236 79704
rect 167288 79750 167362 79778
rect 168116 79784 168190 79812
rect 167460 79756 167512 79762
rect 166816 79620 166868 79626
rect 166816 79562 166868 79568
rect 166722 78840 166778 78849
rect 166722 78775 166778 78784
rect 166552 78628 166672 78656
rect 166552 75954 166580 78628
rect 166828 78305 166856 79562
rect 166908 79484 166960 79490
rect 166908 79426 166960 79432
rect 166920 78713 166948 79426
rect 167000 79416 167052 79422
rect 167000 79358 167052 79364
rect 166906 78704 166962 78713
rect 166906 78639 166962 78648
rect 166814 78296 166870 78305
rect 166814 78231 166870 78240
rect 166632 77308 166684 77314
rect 166632 77250 166684 77256
rect 166540 75948 166592 75954
rect 166540 75890 166592 75896
rect 166540 75404 166592 75410
rect 166540 75346 166592 75352
rect 166448 75336 166500 75342
rect 166448 75278 166500 75284
rect 166276 70366 166396 70394
rect 166172 28620 166224 28626
rect 166172 28562 166224 28568
rect 166080 28484 166132 28490
rect 166080 28426 166132 28432
rect 166276 28422 166304 70366
rect 166552 28830 166580 75346
rect 166644 28898 166672 77250
rect 167012 76022 167040 79358
rect 167000 76016 167052 76022
rect 167000 75958 167052 75964
rect 166724 75948 166776 75954
rect 166724 75890 166776 75896
rect 166632 28892 166684 28898
rect 166632 28834 166684 28840
rect 166540 28824 166592 28830
rect 166540 28766 166592 28772
rect 166264 28416 166316 28422
rect 166264 28358 166316 28364
rect 165896 17400 165948 17406
rect 165896 17342 165948 17348
rect 165804 14544 165856 14550
rect 165804 14486 165856 14492
rect 165712 11824 165764 11830
rect 165712 11766 165764 11772
rect 164240 7608 164292 7614
rect 164240 7550 164292 7556
rect 166078 4856 166134 4865
rect 166078 4791 166134 4800
rect 164882 3496 164938 3505
rect 164882 3431 164938 3440
rect 164896 480 164924 3431
rect 166092 480 166120 4791
rect 166736 3874 166764 75890
rect 167000 75268 167052 75274
rect 167000 75210 167052 75216
rect 167012 58682 167040 75210
rect 167104 68610 167132 79698
rect 167196 78826 167224 79698
rect 167288 79422 167316 79750
rect 167460 79698 167512 79704
rect 167920 79756 167972 79762
rect 167920 79698 167972 79704
rect 167366 79656 167422 79665
rect 167366 79591 167422 79600
rect 167276 79416 167328 79422
rect 167276 79358 167328 79364
rect 167196 78798 167316 78826
rect 167184 78736 167236 78742
rect 167184 78678 167236 78684
rect 167092 68604 167144 68610
rect 167092 68546 167144 68552
rect 167196 68542 167224 78678
rect 167288 72486 167316 78798
rect 167380 78334 167408 79591
rect 167472 78742 167500 79698
rect 167552 79688 167604 79694
rect 167552 79630 167604 79636
rect 167642 79656 167698 79665
rect 167460 78736 167512 78742
rect 167460 78678 167512 78684
rect 167368 78328 167420 78334
rect 167368 78270 167420 78276
rect 167564 78266 167592 79630
rect 167642 79591 167698 79600
rect 167736 79620 167788 79626
rect 167552 78260 167604 78266
rect 167552 78202 167604 78208
rect 167550 78160 167606 78169
rect 167550 78095 167606 78104
rect 167276 72480 167328 72486
rect 167276 72422 167328 72428
rect 167564 71126 167592 78095
rect 167552 71120 167604 71126
rect 167552 71062 167604 71068
rect 167656 70394 167684 79591
rect 167736 79562 167788 79568
rect 167828 79620 167880 79626
rect 167932 79608 167960 79698
rect 168116 79665 168144 79784
rect 168254 79744 168282 80036
rect 168346 79971 168374 80036
rect 168332 79962 168388 79971
rect 168332 79897 168388 79906
rect 168438 79744 168466 80036
rect 168208 79716 168282 79744
rect 168392 79716 168466 79744
rect 168102 79656 168158 79665
rect 167932 79580 168052 79608
rect 168102 79591 168158 79600
rect 167828 79562 167880 79568
rect 167748 71058 167776 79562
rect 167840 75274 167868 79562
rect 168024 77625 168052 79580
rect 168104 79484 168156 79490
rect 168104 79426 168156 79432
rect 168116 79121 168144 79426
rect 168102 79112 168158 79121
rect 168102 79047 168158 79056
rect 168208 78713 168236 79716
rect 168288 79620 168340 79626
rect 168288 79562 168340 79568
rect 168300 78985 168328 79562
rect 168286 78976 168342 78985
rect 168286 78911 168342 78920
rect 168194 78704 168250 78713
rect 168194 78639 168250 78648
rect 168196 77784 168248 77790
rect 168196 77726 168248 77732
rect 168010 77616 168066 77625
rect 168010 77551 168066 77560
rect 168208 77042 168236 77726
rect 168288 77512 168340 77518
rect 168288 77454 168340 77460
rect 168196 77036 168248 77042
rect 168196 76978 168248 76984
rect 168300 75834 168328 77454
rect 168392 77450 168420 79716
rect 168530 79642 168558 80036
rect 168622 79898 168650 80036
rect 168714 79937 168742 80036
rect 168806 79966 168834 80036
rect 168794 79960 168846 79966
rect 168700 79928 168756 79937
rect 168610 79892 168662 79898
rect 168794 79902 168846 79908
rect 168898 79898 168926 80036
rect 168700 79863 168756 79872
rect 168886 79892 168938 79898
rect 168610 79834 168662 79840
rect 168886 79834 168938 79840
rect 168746 79792 168802 79801
rect 168656 79756 168708 79762
rect 168990 79744 169018 80036
rect 168746 79727 168802 79736
rect 168656 79698 168708 79704
rect 168484 79614 168558 79642
rect 168380 77444 168432 77450
rect 168380 77386 168432 77392
rect 168484 76226 168512 79614
rect 168562 79520 168618 79529
rect 168562 79455 168618 79464
rect 168576 79422 168604 79455
rect 168564 79416 168616 79422
rect 168564 79358 168616 79364
rect 168562 79112 168618 79121
rect 168562 79047 168564 79056
rect 168616 79047 168618 79056
rect 168564 79018 168616 79024
rect 168472 76220 168524 76226
rect 168472 76162 168524 76168
rect 168668 76090 168696 79698
rect 168656 76084 168708 76090
rect 168656 76026 168708 76032
rect 168654 75984 168710 75993
rect 168472 75948 168524 75954
rect 168654 75919 168710 75928
rect 168472 75890 168524 75896
rect 168300 75806 168420 75834
rect 167828 75268 167880 75274
rect 167828 75210 167880 75216
rect 168392 72418 168420 75806
rect 168380 72412 168432 72418
rect 168380 72354 168432 72360
rect 167736 71052 167788 71058
rect 167736 70994 167788 71000
rect 167288 70366 167684 70394
rect 167184 68536 167236 68542
rect 167184 68478 167236 68484
rect 167288 68474 167316 70366
rect 167276 68468 167328 68474
rect 167276 68410 167328 68416
rect 167000 58676 167052 58682
rect 167000 58618 167052 58624
rect 168484 8974 168512 75890
rect 168564 74724 168616 74730
rect 168564 74666 168616 74672
rect 168576 20058 168604 74666
rect 168668 20126 168696 75919
rect 168760 29646 168788 79727
rect 168944 79716 169018 79744
rect 169082 79744 169110 80036
rect 169174 79937 169202 80036
rect 169160 79928 169216 79937
rect 169160 79863 169216 79872
rect 169266 79744 169294 80036
rect 169358 79898 169386 80036
rect 169450 79966 169478 80036
rect 169438 79960 169490 79966
rect 169438 79902 169490 79908
rect 169542 79898 169570 80036
rect 169346 79892 169398 79898
rect 169346 79834 169398 79840
rect 169530 79892 169582 79898
rect 169530 79834 169582 79840
rect 169082 79716 169156 79744
rect 168840 79552 168892 79558
rect 168840 79494 168892 79500
rect 168852 60178 168880 79494
rect 168944 75954 168972 79716
rect 169024 79620 169076 79626
rect 169024 79562 169076 79568
rect 168932 75948 168984 75954
rect 168932 75890 168984 75896
rect 169036 73574 169064 79562
rect 169128 75954 169156 79716
rect 169220 79716 169294 79744
rect 169392 79756 169444 79762
rect 169116 75948 169168 75954
rect 169116 75890 169168 75896
rect 169220 75478 169248 79716
rect 169634 79744 169662 80036
rect 169726 79937 169754 80036
rect 169818 79966 169846 80036
rect 169910 79966 169938 80036
rect 170002 79966 170030 80036
rect 170094 79971 170122 80036
rect 169806 79960 169858 79966
rect 169712 79928 169768 79937
rect 169806 79902 169858 79908
rect 169898 79960 169950 79966
rect 169898 79902 169950 79908
rect 169990 79960 170042 79966
rect 169990 79902 170042 79908
rect 170080 79962 170136 79971
rect 170186 79966 170214 80036
rect 170080 79897 170136 79906
rect 170174 79960 170226 79966
rect 170174 79902 170226 79908
rect 169712 79863 169768 79872
rect 170278 79812 170306 80036
rect 170370 79971 170398 80036
rect 170356 79962 170412 79971
rect 170356 79897 170412 79906
rect 170462 79898 170490 80036
rect 170554 79898 170582 80036
rect 170450 79892 170502 79898
rect 170450 79834 170502 79840
rect 170542 79892 170594 79898
rect 170542 79834 170594 79840
rect 170278 79784 170352 79812
rect 169760 79756 169812 79762
rect 169634 79716 169708 79744
rect 169392 79698 169444 79704
rect 169300 79620 169352 79626
rect 169300 79562 169352 79568
rect 169208 75472 169260 75478
rect 169208 75414 169260 75420
rect 169024 73568 169076 73574
rect 169024 73510 169076 73516
rect 169312 70394 169340 79562
rect 169404 75342 169432 79698
rect 169484 79688 169536 79694
rect 169484 79630 169536 79636
rect 169392 75336 169444 75342
rect 169392 75278 169444 75284
rect 169496 74730 169524 79630
rect 169576 79348 169628 79354
rect 169576 79290 169628 79296
rect 169588 79082 169616 79290
rect 169576 79076 169628 79082
rect 169576 79018 169628 79024
rect 169576 78804 169628 78810
rect 169576 78746 169628 78752
rect 169588 77722 169616 78746
rect 169680 78713 169708 79716
rect 169760 79698 169812 79704
rect 170128 79756 170180 79762
rect 170128 79698 170180 79704
rect 169666 78704 169722 78713
rect 169666 78639 169722 78648
rect 169576 77716 169628 77722
rect 169576 77658 169628 77664
rect 169668 75948 169720 75954
rect 169668 75890 169720 75896
rect 169484 74724 169536 74730
rect 169484 74666 169536 74672
rect 169220 70366 169340 70394
rect 169220 68406 169248 70366
rect 169208 68400 169260 68406
rect 169208 68342 169260 68348
rect 168840 60172 168892 60178
rect 168840 60114 168892 60120
rect 168748 29640 168800 29646
rect 168748 29582 168800 29588
rect 168656 20120 168708 20126
rect 168656 20062 168708 20068
rect 168564 20052 168616 20058
rect 168564 19994 168616 20000
rect 168472 8968 168524 8974
rect 168472 8910 168524 8916
rect 169576 5092 169628 5098
rect 169576 5034 169628 5040
rect 166724 3868 166776 3874
rect 166724 3810 166776 3816
rect 167184 3664 167236 3670
rect 167184 3606 167236 3612
rect 167196 480 167224 3606
rect 168378 3360 168434 3369
rect 168378 3295 168434 3304
rect 168392 480 168420 3295
rect 169588 480 169616 5034
rect 169680 4894 169708 75890
rect 169772 10334 169800 79698
rect 170036 79688 170088 79694
rect 169956 79636 170036 79642
rect 169956 79630 170088 79636
rect 169956 79614 170076 79630
rect 169852 76288 169904 76294
rect 169852 76230 169904 76236
rect 169864 11762 169892 76230
rect 169956 21554 169984 79614
rect 170036 79552 170088 79558
rect 170036 79494 170088 79500
rect 169944 21548 169996 21554
rect 169944 21490 169996 21496
rect 170048 21418 170076 79494
rect 170140 79422 170168 79698
rect 170324 79608 170352 79784
rect 170402 79792 170458 79801
rect 170646 79778 170674 80036
rect 170738 79812 170766 80036
rect 170830 79966 170858 80036
rect 170818 79960 170870 79966
rect 170818 79902 170870 79908
rect 170738 79784 170812 79812
rect 170402 79727 170458 79736
rect 170496 79756 170548 79762
rect 170232 79580 170352 79608
rect 170128 79416 170180 79422
rect 170128 79358 170180 79364
rect 170128 78940 170180 78946
rect 170128 78882 170180 78888
rect 170140 78810 170168 78882
rect 170128 78804 170180 78810
rect 170128 78746 170180 78752
rect 170128 78668 170180 78674
rect 170128 78610 170180 78616
rect 170140 78402 170168 78610
rect 170128 78396 170180 78402
rect 170128 78338 170180 78344
rect 170232 76106 170260 79580
rect 170312 79484 170364 79490
rect 170312 79426 170364 79432
rect 170324 78130 170352 79426
rect 170312 78124 170364 78130
rect 170312 78066 170364 78072
rect 170416 77294 170444 79727
rect 170496 79698 170548 79704
rect 170600 79750 170674 79778
rect 170508 79529 170536 79698
rect 170494 79520 170550 79529
rect 170494 79455 170550 79464
rect 170496 79416 170548 79422
rect 170496 79358 170548 79364
rect 170324 77266 170444 77294
rect 170324 76294 170352 77266
rect 170402 77208 170458 77217
rect 170402 77143 170458 77152
rect 170312 76288 170364 76294
rect 170312 76230 170364 76236
rect 170140 76078 170260 76106
rect 170140 21486 170168 76078
rect 170218 75984 170274 75993
rect 170218 75919 170274 75928
rect 170312 75948 170364 75954
rect 170232 25838 170260 75919
rect 170312 75890 170364 75896
rect 170324 68338 170352 75890
rect 170416 69766 170444 77143
rect 170508 73506 170536 79358
rect 170600 75274 170628 79750
rect 170680 79688 170732 79694
rect 170680 79630 170732 79636
rect 170692 77897 170720 79630
rect 170678 77888 170734 77897
rect 170678 77823 170734 77832
rect 170784 75954 170812 79784
rect 170922 79778 170950 80036
rect 171014 79937 171042 80036
rect 171000 79928 171056 79937
rect 171000 79863 171056 79872
rect 170876 79750 170950 79778
rect 170876 75993 170904 79750
rect 171106 79744 171134 80036
rect 171060 79716 171134 79744
rect 171060 78713 171088 79716
rect 171198 79676 171226 80036
rect 171290 79937 171318 80036
rect 171276 79928 171332 79937
rect 171382 79898 171410 80036
rect 171276 79863 171332 79872
rect 171370 79892 171422 79898
rect 171370 79834 171422 79840
rect 171474 79778 171502 80036
rect 171566 79966 171594 80036
rect 171658 79966 171686 80036
rect 171750 79971 171778 80036
rect 171554 79960 171606 79966
rect 171554 79902 171606 79908
rect 171646 79960 171698 79966
rect 171646 79902 171698 79908
rect 171736 79962 171792 79971
rect 171842 79966 171870 80036
rect 171934 79966 171962 80036
rect 172026 79966 172054 80036
rect 171736 79897 171792 79906
rect 171830 79960 171882 79966
rect 171830 79902 171882 79908
rect 171922 79960 171974 79966
rect 171922 79902 171974 79908
rect 172014 79960 172066 79966
rect 172014 79902 172066 79908
rect 172118 79830 172146 80036
rect 172210 79898 172238 80036
rect 172198 79892 172250 79898
rect 172198 79834 172250 79840
rect 172302 79830 172330 80036
rect 172014 79824 172066 79830
rect 172012 79792 172014 79801
rect 172106 79824 172158 79830
rect 172066 79792 172068 79801
rect 171324 79756 171376 79762
rect 171474 79750 171548 79778
rect 171324 79698 171376 79704
rect 171152 79648 171226 79676
rect 171046 78704 171102 78713
rect 171046 78639 171102 78648
rect 171048 78532 171100 78538
rect 171048 78474 171100 78480
rect 170954 78432 171010 78441
rect 170954 78367 171010 78376
rect 170968 77761 170996 78367
rect 170954 77752 171010 77761
rect 170954 77687 171010 77696
rect 171060 77518 171088 78474
rect 171048 77512 171100 77518
rect 171048 77454 171100 77460
rect 170956 76084 171008 76090
rect 170956 76026 171008 76032
rect 170862 75984 170918 75993
rect 170772 75948 170824 75954
rect 170862 75919 170918 75928
rect 170772 75890 170824 75896
rect 170588 75268 170640 75274
rect 170588 75210 170640 75216
rect 170496 73500 170548 73506
rect 170496 73442 170548 73448
rect 170404 69760 170456 69766
rect 170404 69702 170456 69708
rect 170312 68332 170364 68338
rect 170312 68274 170364 68280
rect 170220 25832 170272 25838
rect 170220 25774 170272 25780
rect 170128 21480 170180 21486
rect 170128 21422 170180 21428
rect 170036 21412 170088 21418
rect 170036 21354 170088 21360
rect 170968 20194 170996 76026
rect 171152 75954 171180 79648
rect 171232 79552 171284 79558
rect 171232 79494 171284 79500
rect 171140 75948 171192 75954
rect 171140 75890 171192 75896
rect 171140 75404 171192 75410
rect 171140 75346 171192 75352
rect 170956 20188 171008 20194
rect 170956 20130 171008 20136
rect 169852 11756 169904 11762
rect 169852 11698 169904 11704
rect 169760 10328 169812 10334
rect 169760 10270 169812 10276
rect 169668 4888 169720 4894
rect 169668 4830 169720 4836
rect 171152 4826 171180 75346
rect 171244 17270 171272 79494
rect 171336 17338 171364 79698
rect 171416 79484 171468 79490
rect 171416 79426 171468 79432
rect 171428 19990 171456 79426
rect 171520 78554 171548 79750
rect 171784 79756 171836 79762
rect 172106 79766 172158 79772
rect 172290 79824 172342 79830
rect 172290 79766 172342 79772
rect 172012 79727 172068 79736
rect 172394 79744 172422 80036
rect 172486 79966 172514 80036
rect 172578 79966 172606 80036
rect 172474 79960 172526 79966
rect 172474 79902 172526 79908
rect 172566 79960 172618 79966
rect 172566 79902 172618 79908
rect 172518 79792 172574 79801
rect 172394 79716 172468 79744
rect 172670 79778 172698 80036
rect 172762 79966 172790 80036
rect 172750 79960 172802 79966
rect 172750 79902 172802 79908
rect 172574 79750 172698 79778
rect 172518 79727 172574 79736
rect 171784 79698 171836 79704
rect 171600 79688 171652 79694
rect 171600 79630 171652 79636
rect 171612 78674 171640 79630
rect 171796 79234 171824 79698
rect 172060 79620 172112 79626
rect 172060 79562 172112 79568
rect 171796 79206 171916 79234
rect 171784 79144 171836 79150
rect 171784 79086 171836 79092
rect 171600 78668 171652 78674
rect 171600 78610 171652 78616
rect 171520 78526 171732 78554
rect 171508 78464 171560 78470
rect 171508 78406 171560 78412
rect 171520 77858 171548 78406
rect 171508 77852 171560 77858
rect 171508 77794 171560 77800
rect 171704 76106 171732 78526
rect 171796 78402 171824 79086
rect 171784 78396 171836 78402
rect 171784 78338 171836 78344
rect 171508 76084 171560 76090
rect 171508 76026 171560 76032
rect 171612 76078 171732 76106
rect 171520 25770 171548 76026
rect 171612 28286 171640 76078
rect 171782 75984 171838 75993
rect 171692 75948 171744 75954
rect 171782 75919 171838 75928
rect 171692 75890 171744 75896
rect 171704 28354 171732 75890
rect 171692 28348 171744 28354
rect 171692 28290 171744 28296
rect 171600 28280 171652 28286
rect 171796 28257 171824 75919
rect 171888 60110 171916 79206
rect 172072 75410 172100 79562
rect 172152 79552 172204 79558
rect 172440 79529 172468 79716
rect 172854 79676 172882 80036
rect 172946 79966 172974 80036
rect 172934 79960 172986 79966
rect 172934 79902 172986 79908
rect 173038 79830 173066 80036
rect 173130 79966 173158 80036
rect 173118 79960 173170 79966
rect 173118 79902 173170 79908
rect 173026 79824 173078 79830
rect 173026 79766 173078 79772
rect 172980 79688 173032 79694
rect 172854 79648 172928 79676
rect 172612 79552 172664 79558
rect 172152 79494 172204 79500
rect 172426 79520 172482 79529
rect 172164 78713 172192 79494
rect 172244 79484 172296 79490
rect 172612 79494 172664 79500
rect 172426 79455 172482 79464
rect 172244 79426 172296 79432
rect 172150 78704 172206 78713
rect 172150 78639 172206 78648
rect 172150 78568 172206 78577
rect 172150 78503 172206 78512
rect 172164 76090 172192 78503
rect 172256 76401 172284 79426
rect 172336 79416 172388 79422
rect 172336 79358 172388 79364
rect 172348 78441 172376 79358
rect 172428 79144 172480 79150
rect 172428 79086 172480 79092
rect 172334 78432 172390 78441
rect 172334 78367 172390 78376
rect 172440 77738 172468 79086
rect 172624 78418 172652 79494
rect 172704 79484 172756 79490
rect 172704 79426 172756 79432
rect 172348 77710 172468 77738
rect 172532 78390 172652 78418
rect 172348 77586 172376 77710
rect 172428 77648 172480 77654
rect 172428 77590 172480 77596
rect 172336 77580 172388 77586
rect 172336 77522 172388 77528
rect 172242 76392 172298 76401
rect 172242 76327 172298 76336
rect 172152 76084 172204 76090
rect 172152 76026 172204 76032
rect 172060 75404 172112 75410
rect 172060 75346 172112 75352
rect 172440 70394 172468 77590
rect 172256 70366 172468 70394
rect 172256 64874 172284 70366
rect 171980 64846 172284 64874
rect 171876 60104 171928 60110
rect 171876 60046 171928 60052
rect 171876 58812 171928 58818
rect 171876 58754 171928 58760
rect 171600 28222 171652 28228
rect 171782 28248 171838 28257
rect 171782 28183 171838 28192
rect 171508 25764 171560 25770
rect 171508 25706 171560 25712
rect 171416 19984 171468 19990
rect 171416 19926 171468 19932
rect 171324 17332 171376 17338
rect 171324 17274 171376 17280
rect 171232 17264 171284 17270
rect 171232 17206 171284 17212
rect 170772 4820 170824 4826
rect 170772 4762 170824 4768
rect 171140 4820 171192 4826
rect 171140 4762 171192 4768
rect 170784 480 170812 4762
rect 171888 3262 171916 58754
rect 171980 16574 172008 64846
rect 172532 31278 172560 78390
rect 172612 78192 172664 78198
rect 172612 78134 172664 78140
rect 172520 31272 172572 31278
rect 172520 31214 172572 31220
rect 172624 31210 172652 78134
rect 172716 78062 172744 79426
rect 172796 79416 172848 79422
rect 172796 79358 172848 79364
rect 172704 78056 172756 78062
rect 172704 77998 172756 78004
rect 172808 76634 172836 79358
rect 172900 78946 172928 79648
rect 173222 79642 173250 80036
rect 173314 79898 173342 80036
rect 173406 79937 173434 80036
rect 173498 79966 173526 80036
rect 173590 79966 173618 80036
rect 173682 79966 173710 80036
rect 173774 79971 173802 80036
rect 173486 79960 173538 79966
rect 173392 79928 173448 79937
rect 173302 79892 173354 79898
rect 173486 79902 173538 79908
rect 173578 79960 173630 79966
rect 173578 79902 173630 79908
rect 173670 79960 173722 79966
rect 173670 79902 173722 79908
rect 173760 79962 173816 79971
rect 173866 79966 173894 80036
rect 173760 79897 173816 79906
rect 173854 79960 173906 79966
rect 173854 79902 173906 79908
rect 173392 79863 173448 79872
rect 173302 79834 173354 79840
rect 173578 79824 173630 79830
rect 173958 79812 173986 80036
rect 173912 79784 173986 79812
rect 174050 79812 174078 80036
rect 174142 79971 174170 80036
rect 174128 79962 174184 79971
rect 174234 79966 174262 80036
rect 174326 79966 174354 80036
rect 174418 79966 174446 80036
rect 174510 79966 174538 80036
rect 174602 79966 174630 80036
rect 174128 79897 174184 79906
rect 174222 79960 174274 79966
rect 174222 79902 174274 79908
rect 174314 79960 174366 79966
rect 174314 79902 174366 79908
rect 174406 79960 174458 79966
rect 174406 79902 174458 79908
rect 174498 79960 174550 79966
rect 174498 79902 174550 79908
rect 174590 79960 174642 79966
rect 174694 79937 174722 80036
rect 174786 79966 174814 80036
rect 174878 79966 174906 80036
rect 174774 79960 174826 79966
rect 174590 79902 174642 79908
rect 174680 79928 174736 79937
rect 174774 79902 174826 79908
rect 174866 79960 174918 79966
rect 174970 79937 174998 80036
rect 175062 79966 175090 80036
rect 175050 79960 175102 79966
rect 174866 79902 174918 79908
rect 174956 79928 175012 79937
rect 174680 79863 174736 79872
rect 175050 79902 175102 79908
rect 175154 79898 175182 80036
rect 175246 79971 175274 80036
rect 175232 79962 175288 79971
rect 175338 79966 175366 80036
rect 175430 79971 175458 80036
rect 174956 79863 175012 79872
rect 175142 79892 175194 79898
rect 175232 79897 175288 79906
rect 175326 79960 175378 79966
rect 175326 79902 175378 79908
rect 175416 79962 175472 79971
rect 175416 79897 175472 79906
rect 175142 79834 175194 79840
rect 174774 79824 174826 79830
rect 174050 79784 174124 79812
rect 173630 79772 173848 79778
rect 173578 79766 173848 79772
rect 173590 79750 173848 79766
rect 172980 79630 173032 79636
rect 172888 78940 172940 78946
rect 172888 78882 172940 78888
rect 172888 78532 172940 78538
rect 172888 78474 172940 78480
rect 172796 76628 172848 76634
rect 172796 76570 172848 76576
rect 172704 76424 172756 76430
rect 172704 76366 172756 76372
rect 172612 31204 172664 31210
rect 172612 31146 172664 31152
rect 172716 31142 172744 76366
rect 172796 76356 172848 76362
rect 172796 76298 172848 76304
rect 172704 31136 172756 31142
rect 172704 31078 172756 31084
rect 172808 31074 172836 76298
rect 172900 33862 172928 78474
rect 172992 78198 173020 79630
rect 173176 79614 173250 79642
rect 173532 79688 173584 79694
rect 173532 79630 173584 79636
rect 173624 79688 173676 79694
rect 173624 79630 173676 79636
rect 173440 79620 173492 79626
rect 173176 79422 173204 79614
rect 173440 79562 173492 79568
rect 173256 79552 173308 79558
rect 173256 79494 173308 79500
rect 173346 79520 173402 79529
rect 173164 79416 173216 79422
rect 173164 79358 173216 79364
rect 173072 79348 173124 79354
rect 173072 79290 173124 79296
rect 173084 78606 173112 79290
rect 173164 78940 173216 78946
rect 173164 78882 173216 78888
rect 173072 78600 173124 78606
rect 173072 78542 173124 78548
rect 172980 78192 173032 78198
rect 172980 78134 173032 78140
rect 172980 78056 173032 78062
rect 172980 77998 173032 78004
rect 172992 33930 173020 77998
rect 173176 77294 173204 78882
rect 173268 78656 173296 79494
rect 173346 79455 173402 79464
rect 173360 79286 173388 79455
rect 173348 79280 173400 79286
rect 173348 79222 173400 79228
rect 173268 78628 173388 78656
rect 173176 77266 173296 77294
rect 173072 77172 173124 77178
rect 173072 77114 173124 77120
rect 172980 33924 173032 33930
rect 172980 33866 173032 33872
rect 172888 33856 172940 33862
rect 172888 33798 172940 33804
rect 173084 33794 173112 77114
rect 173164 76628 173216 76634
rect 173164 76570 173216 76576
rect 173176 34066 173204 76570
rect 173164 34060 173216 34066
rect 173164 34002 173216 34008
rect 173268 33998 173296 77266
rect 173360 76430 173388 78628
rect 173452 77994 173480 79562
rect 173440 77988 173492 77994
rect 173440 77930 173492 77936
rect 173348 76424 173400 76430
rect 173348 76366 173400 76372
rect 173544 76362 173572 79630
rect 173636 77178 173664 79630
rect 173716 79552 173768 79558
rect 173716 79494 173768 79500
rect 173728 77353 173756 79494
rect 173820 78538 173848 79750
rect 173808 78532 173860 78538
rect 173808 78474 173860 78480
rect 173808 77444 173860 77450
rect 173808 77386 173860 77392
rect 173714 77344 173770 77353
rect 173714 77279 173770 77288
rect 173624 77172 173676 77178
rect 173624 77114 173676 77120
rect 173532 76356 173584 76362
rect 173532 76298 173584 76304
rect 173820 75478 173848 77386
rect 173808 75472 173860 75478
rect 173808 75414 173860 75420
rect 173912 75138 173940 79784
rect 174096 79642 174124 79784
rect 174772 79792 174774 79801
rect 174826 79792 174828 79801
rect 174452 79756 174504 79762
rect 174372 79716 174452 79744
rect 174096 79614 174216 79642
rect 174084 79552 174136 79558
rect 174084 79494 174136 79500
rect 173992 78056 174044 78062
rect 173992 77998 174044 78004
rect 173900 75132 173952 75138
rect 173900 75074 173952 75080
rect 173256 33992 173308 33998
rect 173256 33934 173308 33940
rect 173072 33788 173124 33794
rect 173072 33730 173124 33736
rect 172796 31068 172848 31074
rect 172796 31010 172848 31016
rect 174004 18630 174032 77998
rect 174096 25634 174124 79494
rect 174188 78577 174216 79614
rect 174174 78568 174230 78577
rect 174174 78503 174230 78512
rect 174266 78432 174322 78441
rect 174266 78367 174322 78376
rect 174174 77888 174230 77897
rect 174174 77823 174230 77832
rect 174188 25702 174216 77823
rect 174176 25696 174228 25702
rect 174176 25638 174228 25644
rect 174084 25628 174136 25634
rect 174084 25570 174136 25576
rect 174280 25566 174308 78367
rect 174372 32434 174400 79716
rect 174772 79727 174828 79736
rect 174910 79792 174966 79801
rect 174910 79727 174966 79736
rect 175096 79756 175148 79762
rect 174452 79698 174504 79704
rect 174544 79620 174596 79626
rect 174596 79580 174676 79608
rect 174544 79562 174596 79568
rect 174452 79552 174504 79558
rect 174452 79494 174504 79500
rect 174464 78062 174492 79494
rect 174544 79484 174596 79490
rect 174544 79426 174596 79432
rect 174452 78056 174504 78062
rect 174452 77998 174504 78004
rect 174452 75132 174504 75138
rect 174452 75074 174504 75080
rect 174464 32502 174492 75074
rect 174556 60042 174584 79426
rect 174648 77897 174676 79580
rect 174728 79552 174780 79558
rect 174728 79494 174780 79500
rect 174634 77888 174690 77897
rect 174634 77823 174690 77832
rect 174740 77772 174768 79494
rect 174820 78668 174872 78674
rect 174820 78610 174872 78616
rect 174648 77744 174768 77772
rect 174648 64190 174676 77744
rect 174832 77654 174860 78610
rect 174820 77648 174872 77654
rect 174820 77590 174872 77596
rect 174924 75914 174952 79727
rect 175096 79698 175148 79704
rect 175188 79756 175240 79762
rect 175522 79744 175550 80036
rect 175188 79698 175240 79704
rect 175476 79716 175550 79744
rect 175004 79280 175056 79286
rect 175004 79222 175056 79228
rect 175016 76537 175044 79222
rect 175002 76528 175058 76537
rect 175002 76463 175058 76472
rect 174740 75886 174952 75914
rect 174740 71774 174768 75886
rect 175108 75313 175136 79698
rect 175200 79121 175228 79698
rect 175372 79688 175424 79694
rect 175372 79630 175424 79636
rect 175280 79144 175332 79150
rect 175186 79112 175242 79121
rect 175280 79086 175332 79092
rect 175186 79047 175242 79056
rect 175186 78704 175242 78713
rect 175186 78639 175242 78648
rect 175094 75304 175150 75313
rect 175094 75239 175150 75248
rect 175096 75200 175148 75206
rect 175096 75142 175148 75148
rect 175108 73030 175136 75142
rect 175096 73024 175148 73030
rect 175096 72966 175148 72972
rect 174740 71746 174860 71774
rect 174636 64184 174688 64190
rect 174636 64126 174688 64132
rect 174544 60036 174596 60042
rect 174544 59978 174596 59984
rect 174452 32496 174504 32502
rect 174452 32438 174504 32444
rect 174360 32428 174412 32434
rect 174360 32370 174412 32376
rect 174268 25560 174320 25566
rect 174268 25502 174320 25508
rect 173992 18624 174044 18630
rect 173992 18566 174044 18572
rect 171980 16546 172100 16574
rect 171968 3528 172020 3534
rect 171968 3470 172020 3476
rect 171876 3256 171928 3262
rect 171876 3198 171928 3204
rect 171980 480 172008 3470
rect 172072 3126 172100 16546
rect 174832 14482 174860 71746
rect 174820 14476 174872 14482
rect 174820 14418 174872 14424
rect 175200 6254 175228 78639
rect 175292 77178 175320 79086
rect 175384 78198 175412 79630
rect 175476 79506 175504 79716
rect 175614 79676 175642 80036
rect 175706 79812 175734 80036
rect 175798 79971 175826 80036
rect 175784 79962 175840 79971
rect 175784 79897 175840 79906
rect 175706 79784 175780 79812
rect 175614 79648 175688 79676
rect 175476 79478 175596 79506
rect 175464 79416 175516 79422
rect 175464 79358 175516 79364
rect 175372 78192 175424 78198
rect 175372 78134 175424 78140
rect 175476 77704 175504 79358
rect 175568 78441 175596 79478
rect 175660 78538 175688 79648
rect 175648 78532 175700 78538
rect 175648 78474 175700 78480
rect 175554 78432 175610 78441
rect 175554 78367 175610 78376
rect 175752 78130 175780 79784
rect 175890 79744 175918 80036
rect 175982 79966 176010 80036
rect 175970 79960 176022 79966
rect 175970 79902 176022 79908
rect 176074 79898 176102 80036
rect 176166 79966 176194 80036
rect 176154 79960 176206 79966
rect 176154 79902 176206 79908
rect 176062 79892 176114 79898
rect 176062 79834 176114 79840
rect 175844 79716 175918 79744
rect 176016 79756 176068 79762
rect 175844 78674 175872 79716
rect 176016 79698 176068 79704
rect 176108 79756 176160 79762
rect 176258 79744 176286 80036
rect 176350 79966 176378 80036
rect 176338 79960 176390 79966
rect 176442 79937 176470 80036
rect 176534 79966 176562 80036
rect 176626 79966 176654 80036
rect 176718 79966 176746 80036
rect 176810 79966 176838 80036
rect 176902 79966 176930 80036
rect 176994 79966 177022 80036
rect 177086 79966 177114 80036
rect 176522 79960 176574 79966
rect 176338 79902 176390 79908
rect 176428 79928 176484 79937
rect 176522 79902 176574 79908
rect 176614 79960 176666 79966
rect 176614 79902 176666 79908
rect 176706 79960 176758 79966
rect 176706 79902 176758 79908
rect 176798 79960 176850 79966
rect 176798 79902 176850 79908
rect 176890 79960 176942 79966
rect 176890 79902 176942 79908
rect 176982 79960 177034 79966
rect 176982 79902 177034 79908
rect 177074 79960 177126 79966
rect 177178 79937 177206 80036
rect 177270 79966 177298 80036
rect 177362 79966 177390 80036
rect 177258 79960 177310 79966
rect 177074 79902 177126 79908
rect 177164 79928 177220 79937
rect 176428 79863 176484 79872
rect 177258 79902 177310 79908
rect 177350 79960 177402 79966
rect 177350 79902 177402 79908
rect 177454 79898 177482 80036
rect 177164 79863 177220 79872
rect 177442 79892 177494 79898
rect 177442 79834 177494 79840
rect 177304 79824 177356 79830
rect 177118 79792 177174 79801
rect 176108 79698 176160 79704
rect 176212 79716 176286 79744
rect 176476 79756 176528 79762
rect 176028 78713 176056 79698
rect 176014 78704 176070 78713
rect 175832 78668 175884 78674
rect 176014 78639 176070 78648
rect 175832 78610 175884 78616
rect 175740 78124 175792 78130
rect 175740 78066 175792 78072
rect 175832 78056 175884 78062
rect 175832 77998 175884 78004
rect 175384 77676 175504 77704
rect 175280 77172 175332 77178
rect 175280 77114 175332 77120
rect 175384 75313 175412 77676
rect 175648 76220 175700 76226
rect 175648 76162 175700 76168
rect 175462 75984 175518 75993
rect 175462 75919 175518 75928
rect 175370 75304 175426 75313
rect 175370 75239 175426 75248
rect 175476 70394 175504 75919
rect 175660 70394 175688 76162
rect 175292 70366 175504 70394
rect 175568 70366 175688 70394
rect 175844 70394 175872 77998
rect 175924 77988 175976 77994
rect 175924 77930 175976 77936
rect 175936 75206 175964 77930
rect 176016 76016 176068 76022
rect 176016 75958 176068 75964
rect 175924 75200 175976 75206
rect 175924 75142 175976 75148
rect 176028 70394 176056 75958
rect 176120 73166 176148 79698
rect 176212 79014 176240 79716
rect 176476 79698 176528 79704
rect 176568 79756 176620 79762
rect 176568 79698 176620 79704
rect 176844 79756 176896 79762
rect 176844 79698 176896 79704
rect 176936 79756 176988 79762
rect 176988 79716 177068 79744
rect 177546 79778 177574 80036
rect 177304 79766 177356 79772
rect 177118 79727 177174 79736
rect 177212 79756 177264 79762
rect 176936 79698 176988 79704
rect 176384 79688 176436 79694
rect 176384 79630 176436 79636
rect 176396 79286 176424 79630
rect 176384 79280 176436 79286
rect 176384 79222 176436 79228
rect 176292 79212 176344 79218
rect 176292 79154 176344 79160
rect 176200 79008 176252 79014
rect 176200 78950 176252 78956
rect 176200 77920 176252 77926
rect 176200 77862 176252 77868
rect 176212 76650 176240 77862
rect 176304 76809 176332 79154
rect 176488 77994 176516 79698
rect 176580 78713 176608 79698
rect 176856 79642 176884 79698
rect 176856 79614 176976 79642
rect 176844 79552 176896 79558
rect 176844 79494 176896 79500
rect 176752 79348 176804 79354
rect 176752 79290 176804 79296
rect 176660 79076 176712 79082
rect 176660 79018 176712 79024
rect 176672 78849 176700 79018
rect 176658 78840 176714 78849
rect 176658 78775 176714 78784
rect 176566 78704 176622 78713
rect 176566 78639 176622 78648
rect 176764 78538 176792 79290
rect 176568 78532 176620 78538
rect 176568 78474 176620 78480
rect 176752 78532 176804 78538
rect 176752 78474 176804 78480
rect 176476 77988 176528 77994
rect 176476 77930 176528 77936
rect 176384 77784 176436 77790
rect 176384 77726 176436 77732
rect 176474 77752 176530 77761
rect 176290 76800 176346 76809
rect 176290 76735 176346 76744
rect 176212 76622 176332 76650
rect 176200 75676 176252 75682
rect 176200 75618 176252 75624
rect 176108 73160 176160 73166
rect 176108 73102 176160 73108
rect 175844 70366 175964 70394
rect 176028 70366 176148 70394
rect 175292 44878 175320 70366
rect 175280 44872 175332 44878
rect 175280 44814 175332 44820
rect 175188 6248 175240 6254
rect 175188 6190 175240 6196
rect 173164 5024 173216 5030
rect 173164 4966 173216 4972
rect 172060 3120 172112 3126
rect 172060 3062 172112 3068
rect 173176 480 173204 4966
rect 174268 3596 174320 3602
rect 174268 3538 174320 3544
rect 174280 480 174308 3538
rect 175464 3460 175516 3466
rect 175464 3402 175516 3408
rect 175476 480 175504 3402
rect 175568 3058 175596 70366
rect 175936 3330 175964 70366
rect 176120 3806 176148 70366
rect 176108 3800 176160 3806
rect 176108 3742 176160 3748
rect 176212 3534 176240 75618
rect 176304 15910 176332 76622
rect 176396 36582 176424 77726
rect 176474 77687 176530 77696
rect 176488 77489 176516 77687
rect 176474 77480 176530 77489
rect 176474 77415 176530 77424
rect 176474 73536 176530 73545
rect 176474 73471 176530 73480
rect 176488 69698 176516 73471
rect 176476 69692 176528 69698
rect 176476 69634 176528 69640
rect 176384 36576 176436 36582
rect 176384 36518 176436 36524
rect 176292 15904 176344 15910
rect 176292 15846 176344 15852
rect 176580 6186 176608 78474
rect 176856 77353 176884 79494
rect 176948 78849 176976 79614
rect 176934 78840 176990 78849
rect 176934 78775 176990 78784
rect 177040 78305 177068 79716
rect 177132 79354 177160 79727
rect 177212 79698 177264 79704
rect 177224 79393 177252 79698
rect 177210 79384 177266 79393
rect 177120 79348 177172 79354
rect 177210 79319 177266 79328
rect 177120 79290 177172 79296
rect 177316 79218 177344 79766
rect 177500 79750 177574 79778
rect 177396 79484 177448 79490
rect 177396 79426 177448 79432
rect 177304 79212 177356 79218
rect 177304 79154 177356 79160
rect 177118 79112 177174 79121
rect 177118 79047 177174 79056
rect 177026 78296 177082 78305
rect 177026 78231 177082 78240
rect 177132 78169 177160 79047
rect 177408 78674 177436 79426
rect 177500 79121 177528 79750
rect 177638 79744 177666 80036
rect 177730 79898 177758 80036
rect 177718 79892 177770 79898
rect 177718 79834 177770 79840
rect 177822 79830 177850 80036
rect 177810 79824 177862 79830
rect 177914 79812 177942 80036
rect 178006 79937 178034 80036
rect 177992 79928 178048 79937
rect 177992 79863 178048 79872
rect 177914 79801 177988 79812
rect 177914 79792 178002 79801
rect 177914 79784 177946 79792
rect 177810 79766 177862 79772
rect 177638 79716 177712 79744
rect 178098 79744 178126 80036
rect 177946 79727 178002 79736
rect 177684 79529 177712 79716
rect 178052 79716 178126 79744
rect 178052 79665 178080 79716
rect 178190 79676 178218 80036
rect 178282 79744 178310 80036
rect 178374 79812 178402 80036
rect 178466 79966 178494 80036
rect 178454 79960 178506 79966
rect 178558 79937 178586 80036
rect 178454 79902 178506 79908
rect 178544 79928 178600 79937
rect 178544 79863 178600 79872
rect 178374 79784 178540 79812
rect 178282 79716 178356 79744
rect 178038 79656 178094 79665
rect 178190 79648 178264 79676
rect 178038 79591 178094 79600
rect 177670 79520 177726 79529
rect 177670 79455 177726 79464
rect 178040 79484 178092 79490
rect 178040 79426 178092 79432
rect 178132 79484 178184 79490
rect 178132 79426 178184 79432
rect 177486 79112 177542 79121
rect 177486 79047 177542 79056
rect 178052 78878 178080 79426
rect 178144 79082 178172 79426
rect 178236 79257 178264 79648
rect 178222 79248 178278 79257
rect 178222 79183 178278 79192
rect 178132 79076 178184 79082
rect 178132 79018 178184 79024
rect 177856 78872 177908 78878
rect 177856 78814 177908 78820
rect 178040 78872 178092 78878
rect 178040 78814 178092 78820
rect 177764 78736 177816 78742
rect 177764 78678 177816 78684
rect 177212 78668 177264 78674
rect 177212 78610 177264 78616
rect 177396 78668 177448 78674
rect 177396 78610 177448 78616
rect 177118 78160 177174 78169
rect 177118 78095 177174 78104
rect 177224 77926 177252 78610
rect 177212 77920 177264 77926
rect 177212 77862 177264 77868
rect 177304 77852 177356 77858
rect 177304 77794 177356 77800
rect 177212 77716 177264 77722
rect 177212 77658 177264 77664
rect 176842 77344 176898 77353
rect 176842 77279 176898 77288
rect 177224 49026 177252 77658
rect 177316 73846 177344 77794
rect 177578 77752 177634 77761
rect 177578 77687 177634 77696
rect 177488 77512 177540 77518
rect 177488 77454 177540 77460
rect 177394 75848 177450 75857
rect 177394 75783 177450 75792
rect 177304 73840 177356 73846
rect 177304 73782 177356 73788
rect 177304 73568 177356 73574
rect 177304 73510 177356 73516
rect 177212 49020 177264 49026
rect 177212 48962 177264 48968
rect 176568 6180 176620 6186
rect 176568 6122 176620 6128
rect 177316 3602 177344 73510
rect 177408 3670 177436 75783
rect 177500 9246 177528 77454
rect 177488 9240 177540 9246
rect 177488 9182 177540 9188
rect 177592 3738 177620 77687
rect 177672 77376 177724 77382
rect 177672 77318 177724 77324
rect 177684 74610 177712 77318
rect 177776 75682 177804 78678
rect 177868 76634 177896 78814
rect 178328 78169 178356 79716
rect 178406 79248 178462 79257
rect 178406 79183 178462 79192
rect 178420 78810 178448 79183
rect 178512 78985 178540 79784
rect 178650 79642 178678 80036
rect 178742 79744 178770 80036
rect 178834 79812 178862 80036
rect 178926 79966 178954 80036
rect 178914 79960 178966 79966
rect 178914 79902 178966 79908
rect 178834 79784 178908 79812
rect 178742 79716 178816 79744
rect 178604 79614 178678 79642
rect 178498 78976 178554 78985
rect 178604 78946 178632 79614
rect 178498 78911 178554 78920
rect 178592 78940 178644 78946
rect 178592 78882 178644 78888
rect 178408 78804 178460 78810
rect 178408 78746 178460 78752
rect 178788 78606 178816 79716
rect 178880 79150 178908 79784
rect 179018 79778 179046 80036
rect 179110 79971 179138 80036
rect 179096 79962 179152 79971
rect 179096 79897 179152 79906
rect 179018 79750 179092 79778
rect 178868 79144 178920 79150
rect 178868 79086 178920 79092
rect 178776 78600 178828 78606
rect 178776 78542 178828 78548
rect 178314 78160 178370 78169
rect 178314 78095 178370 78104
rect 178038 78024 178094 78033
rect 178038 77959 178094 77968
rect 178052 77466 178080 77959
rect 178776 77648 178828 77654
rect 178776 77590 178828 77596
rect 177960 77438 178080 77466
rect 177856 76628 177908 76634
rect 177856 76570 177908 76576
rect 177764 75676 177816 75682
rect 177764 75618 177816 75624
rect 177684 74582 177896 74610
rect 177672 73840 177724 73846
rect 177672 73782 177724 73788
rect 177684 21622 177712 73782
rect 177764 73500 177816 73506
rect 177764 73442 177816 73448
rect 177672 21616 177724 21622
rect 177672 21558 177724 21564
rect 177580 3732 177632 3738
rect 177580 3674 177632 3680
rect 177396 3664 177448 3670
rect 177396 3606 177448 3612
rect 177304 3596 177356 3602
rect 177304 3538 177356 3544
rect 176200 3528 176252 3534
rect 176200 3470 176252 3476
rect 177776 3466 177804 73442
rect 177868 39370 177896 74582
rect 177960 43450 177988 77438
rect 178224 77308 178276 77314
rect 178224 77250 178276 77256
rect 178132 75064 178184 75070
rect 178132 75006 178184 75012
rect 178040 73636 178092 73642
rect 178040 73578 178092 73584
rect 178052 70378 178080 73578
rect 178040 70372 178092 70378
rect 178040 70314 178092 70320
rect 178040 69624 178092 69630
rect 178040 69566 178092 69572
rect 177948 43444 178000 43450
rect 177948 43386 178000 43392
rect 177856 39364 177908 39370
rect 177856 39306 177908 39312
rect 178052 16574 178080 69566
rect 178144 22914 178172 75006
rect 178236 45558 178264 77250
rect 178500 76492 178552 76498
rect 178500 76434 178552 76440
rect 178512 72350 178540 76434
rect 178788 73846 178816 77590
rect 179064 77489 179092 79750
rect 179202 79744 179230 80036
rect 179294 79898 179322 80036
rect 179282 79892 179334 79898
rect 179282 79834 179334 79840
rect 179386 79778 179414 80036
rect 179972 80028 180024 80034
rect 179972 79970 180024 79976
rect 179696 79960 179748 79966
rect 179696 79902 179748 79908
rect 179156 79716 179230 79744
rect 179340 79750 179414 79778
rect 179156 78538 179184 79716
rect 179340 79642 179368 79750
rect 179248 79614 179368 79642
rect 179144 78532 179196 78538
rect 179144 78474 179196 78480
rect 179050 77480 179106 77489
rect 179050 77415 179106 77424
rect 179144 76288 179196 76294
rect 179144 76230 179196 76236
rect 179052 76152 179104 76158
rect 179052 76094 179104 76100
rect 178958 74896 179014 74905
rect 178958 74831 179014 74840
rect 178866 74216 178922 74225
rect 178866 74151 178922 74160
rect 178776 73840 178828 73846
rect 178776 73782 178828 73788
rect 178500 72344 178552 72350
rect 178500 72286 178552 72292
rect 178316 71256 178368 71262
rect 178316 71198 178368 71204
rect 178328 69630 178356 71198
rect 178880 69630 178908 74151
rect 178316 69624 178368 69630
rect 178316 69566 178368 69572
rect 178868 69624 178920 69630
rect 178868 69566 178920 69572
rect 178972 68746 179000 74831
rect 179064 71262 179092 76094
rect 179156 71670 179184 76230
rect 179248 75070 179276 79614
rect 179708 78441 179736 79902
rect 179788 79892 179840 79898
rect 179788 79834 179840 79840
rect 179694 78432 179750 78441
rect 179694 78367 179750 78376
rect 179800 77314 179828 79834
rect 179984 79354 180012 79970
rect 180248 79824 180300 79830
rect 180248 79766 180300 79772
rect 180614 79792 180670 79801
rect 179972 79348 180024 79354
rect 179972 79290 180024 79296
rect 179880 79280 179932 79286
rect 179880 79222 179932 79228
rect 179892 79082 179920 79222
rect 179880 79076 179932 79082
rect 179880 79018 179932 79024
rect 179878 78568 179934 78577
rect 180260 78538 180288 79766
rect 180524 79756 180576 79762
rect 180614 79727 180670 79736
rect 180524 79698 180576 79704
rect 180536 79286 180564 79698
rect 180524 79280 180576 79286
rect 180524 79222 180576 79228
rect 180522 78976 180578 78985
rect 180522 78911 180578 78920
rect 180536 78878 180564 78911
rect 180524 78872 180576 78878
rect 180524 78814 180576 78820
rect 179878 78503 179934 78512
rect 180248 78532 180300 78538
rect 179892 78198 179920 78503
rect 180248 78474 180300 78480
rect 179880 78192 179932 78198
rect 179880 78134 179932 78140
rect 180628 77586 180656 79727
rect 181720 79620 181772 79626
rect 181720 79562 181772 79568
rect 181732 79218 181760 79562
rect 181720 79212 181772 79218
rect 181720 79154 181772 79160
rect 188908 78538 188936 80038
rect 188896 78532 188948 78538
rect 188896 78474 188948 78480
rect 189000 78305 189028 80650
rect 188986 78296 189042 78305
rect 188986 78231 189042 78240
rect 187884 77988 187936 77994
rect 187884 77930 187936 77936
rect 187896 77858 187924 77930
rect 187884 77852 187936 77858
rect 187884 77794 187936 77800
rect 180616 77580 180668 77586
rect 180616 77522 180668 77528
rect 189092 77353 189120 80718
rect 189078 77344 189134 77353
rect 179788 77308 179840 77314
rect 189078 77279 189134 77288
rect 179788 77250 179840 77256
rect 185032 77240 185084 77246
rect 185032 77182 185084 77188
rect 181442 76664 181498 76673
rect 181442 76599 181498 76608
rect 181456 76401 181484 76599
rect 181442 76392 181498 76401
rect 181442 76327 181498 76336
rect 179236 75064 179288 75070
rect 179236 75006 179288 75012
rect 179418 75032 179474 75041
rect 179418 74967 179474 74976
rect 179144 71664 179196 71670
rect 179144 71606 179196 71612
rect 179052 71256 179104 71262
rect 179052 71198 179104 71204
rect 179432 69562 179460 74967
rect 179420 69556 179472 69562
rect 179420 69498 179472 69504
rect 181996 69488 182048 69494
rect 181996 69430 182048 69436
rect 178960 68740 179012 68746
rect 178960 68682 179012 68688
rect 179418 68504 179474 68513
rect 179418 68439 179474 68448
rect 178224 45552 178276 45558
rect 178224 45494 178276 45500
rect 178132 22908 178184 22914
rect 178132 22850 178184 22856
rect 179432 16574 179460 68439
rect 182008 67114 182036 69430
rect 181996 67108 182048 67114
rect 181996 67050 182048 67056
rect 182178 66872 182234 66881
rect 182178 66807 182234 66816
rect 178052 16546 178632 16574
rect 179432 16546 180288 16574
rect 177856 3528 177908 3534
rect 177856 3470 177908 3476
rect 177948 3528 178000 3534
rect 177948 3470 178000 3476
rect 177764 3460 177816 3466
rect 177764 3402 177816 3408
rect 175924 3324 175976 3330
rect 175924 3266 175976 3272
rect 176660 3256 176712 3262
rect 176660 3198 176712 3204
rect 175556 3052 175608 3058
rect 175556 2994 175608 3000
rect 176672 480 176700 3198
rect 177868 480 177896 3470
rect 177960 3330 177988 3470
rect 177948 3324 178000 3330
rect 177948 3266 178000 3272
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 180260 480 180288 16546
rect 181444 3664 181496 3670
rect 181444 3606 181496 3612
rect 181456 480 181484 3606
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182192 354 182220 66807
rect 183558 57216 183614 57225
rect 183558 57151 183614 57160
rect 183572 16574 183600 57151
rect 183572 16546 183784 16574
rect 183756 480 183784 16546
rect 185044 6914 185072 77182
rect 187700 32700 187752 32706
rect 187700 32642 187752 32648
rect 186320 26104 186372 26110
rect 186320 26046 186372 26052
rect 186332 16574 186360 26046
rect 187712 16574 187740 32642
rect 189184 24138 189212 129746
rect 189276 126954 189304 201486
rect 189356 160744 189408 160750
rect 189356 160686 189408 160692
rect 189264 126948 189316 126954
rect 189264 126890 189316 126896
rect 189368 122834 189396 160686
rect 189448 145580 189500 145586
rect 189448 145522 189500 145528
rect 189276 122806 189396 122834
rect 189276 116634 189304 122806
rect 189356 121440 189408 121446
rect 189356 121382 189408 121388
rect 189368 120737 189396 121382
rect 189354 120728 189410 120737
rect 189354 120663 189410 120672
rect 189354 116648 189410 116657
rect 189276 116606 189354 116634
rect 189354 116583 189410 116592
rect 189460 113937 189488 145522
rect 189540 144288 189592 144294
rect 189540 144230 189592 144236
rect 189446 113928 189502 113937
rect 189446 113863 189502 113872
rect 189552 112577 189580 144230
rect 189630 130520 189686 130529
rect 189630 130455 189686 130464
rect 189644 129810 189672 130455
rect 189632 129804 189684 129810
rect 189632 129746 189684 129752
rect 189632 126948 189684 126954
rect 189632 126890 189684 126896
rect 189644 126177 189672 126890
rect 189630 126168 189686 126177
rect 189630 126103 189686 126112
rect 189736 119377 189764 462334
rect 189722 119368 189778 119377
rect 189722 119303 189778 119312
rect 189538 112568 189594 112577
rect 189538 112503 189594 112512
rect 189724 111852 189776 111858
rect 189724 111794 189776 111800
rect 189354 82376 189410 82385
rect 189354 82311 189410 82320
rect 189368 77625 189396 82311
rect 189736 79422 189764 111794
rect 189724 79416 189776 79422
rect 189724 79358 189776 79364
rect 189354 77616 189410 77625
rect 190472 77586 190500 700266
rect 190552 514820 190604 514826
rect 190552 514762 190604 514768
rect 190564 117473 190592 514762
rect 190644 253972 190696 253978
rect 190644 253914 190696 253920
rect 190656 124273 190684 253914
rect 191196 148368 191248 148374
rect 191196 148310 191248 148316
rect 190828 146940 190880 146946
rect 190828 146882 190880 146888
rect 190734 129704 190790 129713
rect 190734 129639 190790 129648
rect 190642 124264 190698 124273
rect 190642 124199 190698 124208
rect 190550 117464 190606 117473
rect 190550 117399 190606 117408
rect 189354 77551 189410 77560
rect 190460 77580 190512 77586
rect 190460 77522 190512 77528
rect 190748 69902 190776 129639
rect 190840 114753 190868 146882
rect 191104 142928 191156 142934
rect 191104 142870 191156 142876
rect 191012 141500 191064 141506
rect 191012 141442 191064 141448
rect 190920 140208 190972 140214
rect 190920 140150 190972 140156
rect 190826 114744 190882 114753
rect 190826 114679 190882 114688
rect 190932 109313 190960 140150
rect 191024 110673 191052 141442
rect 191116 121553 191144 142870
rect 191208 126993 191236 148310
rect 192024 140548 192076 140554
rect 192024 140490 192076 140496
rect 191932 139460 191984 139466
rect 191932 139402 191984 139408
rect 191944 128353 191972 139402
rect 191930 128344 191986 128353
rect 191930 128279 191986 128288
rect 191194 126984 191250 126993
rect 191194 126919 191250 126928
rect 192036 122913 192064 140490
rect 192022 122904 192078 122913
rect 192022 122839 192078 122848
rect 191102 121544 191158 121553
rect 191102 121479 191158 121488
rect 191010 110664 191066 110673
rect 191010 110599 191066 110608
rect 190918 109304 190974 109313
rect 190918 109239 190974 109248
rect 191932 108996 191984 109002
rect 191932 108938 191984 108944
rect 191944 107953 191972 108938
rect 191930 107944 191986 107953
rect 191930 107879 191986 107888
rect 191932 107636 191984 107642
rect 191932 107578 191984 107584
rect 191944 106593 191972 107578
rect 191930 106584 191986 106593
rect 191930 106519 191986 106528
rect 191932 106276 191984 106282
rect 191932 106218 191984 106224
rect 191944 105233 191972 106218
rect 191930 105224 191986 105233
rect 191930 105159 191986 105168
rect 191932 101176 191984 101182
rect 191930 101144 191932 101153
rect 191984 101144 191986 101153
rect 191930 101079 191986 101088
rect 192392 100700 192444 100706
rect 192392 100642 192444 100648
rect 192404 99793 192432 100642
rect 192390 99784 192446 99793
rect 192390 99719 192446 99728
rect 192116 98524 192168 98530
rect 192116 98466 192168 98472
rect 192128 98433 192156 98466
rect 192114 98424 192170 98433
rect 192114 98359 192170 98368
rect 192208 97504 192260 97510
rect 192208 97446 192260 97452
rect 192220 97073 192248 97446
rect 192206 97064 192262 97073
rect 192206 96999 192262 97008
rect 191932 96484 191984 96490
rect 191932 96426 191984 96432
rect 191944 95713 191972 96426
rect 191930 95704 191986 95713
rect 191930 95639 191986 95648
rect 192496 79286 192524 700606
rect 200764 700460 200816 700466
rect 200764 700402 200816 700408
rect 199384 700392 199436 700398
rect 199384 700334 199436 700340
rect 198004 700324 198056 700330
rect 198004 700266 198056 700272
rect 193864 699712 193916 699718
rect 193864 699654 193916 699660
rect 192576 418192 192628 418198
rect 192576 418134 192628 418140
rect 192588 92993 192616 418134
rect 192668 191888 192720 191894
rect 192668 191830 192720 191836
rect 192574 92984 192630 92993
rect 192574 92919 192630 92928
rect 192574 82104 192630 82113
rect 192574 82039 192630 82048
rect 192484 79280 192536 79286
rect 192484 79222 192536 79228
rect 191840 75812 191892 75818
rect 191840 75754 191892 75760
rect 190736 69896 190788 69902
rect 190736 69838 190788 69844
rect 189172 24132 189224 24138
rect 189172 24074 189224 24080
rect 191852 16574 191880 75754
rect 192588 60722 192616 82039
rect 192680 79150 192708 191830
rect 192760 151836 192812 151842
rect 192760 151778 192812 151784
rect 192668 79144 192720 79150
rect 192668 79086 192720 79092
rect 192772 79014 192800 151778
rect 193128 104848 193180 104854
rect 193128 104790 193180 104796
rect 193140 103873 193168 104790
rect 193126 103864 193182 103873
rect 193126 103799 193182 103808
rect 193128 102536 193180 102542
rect 193126 102504 193128 102513
rect 193180 102504 193182 102513
rect 193126 102439 193182 102448
rect 193128 95192 193180 95198
rect 193128 95134 193180 95140
rect 193140 94353 193168 95134
rect 193126 94344 193182 94353
rect 193126 94279 193182 94288
rect 193128 92472 193180 92478
rect 193128 92414 193180 92420
rect 193140 91633 193168 92414
rect 193126 91624 193182 91633
rect 193126 91559 193182 91568
rect 193128 91044 193180 91050
rect 193128 90986 193180 90992
rect 193140 90273 193168 90986
rect 193126 90264 193182 90273
rect 193126 90199 193182 90208
rect 193128 89684 193180 89690
rect 193128 89626 193180 89632
rect 192944 89004 192996 89010
rect 192944 88946 192996 88952
rect 192956 87553 192984 88946
rect 193140 88913 193168 89626
rect 193126 88904 193182 88913
rect 193126 88839 193182 88848
rect 193036 87644 193088 87650
rect 193036 87586 193088 87592
rect 192942 87544 192998 87553
rect 192942 87479 192998 87488
rect 193048 86193 193076 87586
rect 193034 86184 193090 86193
rect 193034 86119 193090 86128
rect 193128 85536 193180 85542
rect 193128 85478 193180 85484
rect 193140 84833 193168 85478
rect 193126 84824 193182 84833
rect 193126 84759 193182 84768
rect 193128 84176 193180 84182
rect 193128 84118 193180 84124
rect 193140 83473 193168 84118
rect 193126 83464 193182 83473
rect 193126 83399 193182 83408
rect 193126 80744 193182 80753
rect 193126 80679 193182 80688
rect 193140 80170 193168 80679
rect 193128 80164 193180 80170
rect 193128 80106 193180 80112
rect 193876 79218 193904 699654
rect 196624 683188 196676 683194
rect 196624 683130 196676 683136
rect 193956 630692 194008 630698
rect 193956 630634 194008 630640
rect 193968 98530 193996 630634
rect 194048 576904 194100 576910
rect 194048 576846 194100 576852
rect 193956 98524 194008 98530
rect 193956 98466 194008 98472
rect 194060 97510 194088 576846
rect 194140 524476 194192 524482
rect 194140 524418 194192 524424
rect 194048 97504 194100 97510
rect 194048 97446 194100 97452
rect 194152 96490 194180 524418
rect 194232 231872 194284 231878
rect 194232 231814 194284 231820
rect 194140 96484 194192 96490
rect 194140 96426 194192 96432
rect 194244 79830 194272 231814
rect 196636 100706 196664 683130
rect 198016 101182 198044 700266
rect 199396 102542 199424 700334
rect 200776 104854 200804 700402
rect 202800 699718 202828 703520
rect 218992 700738 219020 703520
rect 207664 700732 207716 700738
rect 207664 700674 207716 700680
rect 218980 700732 219032 700738
rect 218980 700674 219032 700680
rect 206284 700596 206336 700602
rect 206284 700538 206336 700544
rect 203524 700528 203576 700534
rect 203524 700470 203576 700476
rect 202788 699712 202840 699718
rect 202788 699654 202840 699660
rect 202144 258120 202196 258126
rect 202144 258062 202196 258068
rect 200764 104848 200816 104854
rect 200764 104790 200816 104796
rect 199384 102536 199436 102542
rect 199384 102478 199436 102484
rect 198004 101176 198056 101182
rect 198004 101118 198056 101124
rect 196624 100700 196676 100706
rect 196624 100642 196676 100648
rect 202156 89690 202184 258062
rect 203536 106282 203564 700470
rect 206296 107642 206324 700538
rect 207676 109002 207704 700674
rect 221464 470620 221516 470626
rect 221464 470562 221516 470568
rect 207664 108996 207716 109002
rect 207664 108938 207716 108944
rect 206284 107636 206336 107642
rect 206284 107578 206336 107584
rect 203524 106276 203576 106282
rect 203524 106218 203576 106224
rect 221476 95198 221504 470562
rect 225604 218068 225656 218074
rect 225604 218010 225656 218016
rect 224224 178084 224276 178090
rect 224224 178026 224276 178032
rect 221464 95192 221516 95198
rect 221464 95134 221516 95140
rect 202144 89684 202196 89690
rect 202144 89626 202196 89632
rect 224236 87650 224264 178026
rect 225616 89010 225644 218010
rect 234632 147014 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700670 267688 703520
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 234620 147008 234672 147014
rect 234620 146950 234672 146956
rect 299492 145654 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 299480 145648 299532 145654
rect 299480 145590 299532 145596
rect 225604 89004 225656 89010
rect 225604 88946 225656 88952
rect 224224 87644 224276 87650
rect 224224 87586 224276 87592
rect 194232 79824 194284 79830
rect 194232 79766 194284 79772
rect 331232 79529 331260 702986
rect 348804 700534 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 360844 364404 360896 364410
rect 360844 364346 360896 364352
rect 359464 311908 359516 311914
rect 359464 311850 359516 311856
rect 359476 91050 359504 311850
rect 359556 94512 359608 94518
rect 359556 94454 359608 94460
rect 359464 91044 359516 91050
rect 359464 90986 359516 90992
rect 359568 84182 359596 94454
rect 360856 92478 360884 364346
rect 364352 144226 364380 702406
rect 364340 144220 364392 144226
rect 364340 144162 364392 144168
rect 360936 94580 360988 94586
rect 360936 94522 360988 94528
rect 360844 92472 360896 92478
rect 360844 92414 360896 92420
rect 360948 85542 360976 94522
rect 360936 85536 360988 85542
rect 360936 85478 360988 85484
rect 359556 84176 359608 84182
rect 359556 84118 359608 84124
rect 331218 79520 331274 79529
rect 331218 79455 331274 79464
rect 193864 79212 193916 79218
rect 193864 79154 193916 79160
rect 397472 79121 397500 703520
rect 413664 700466 413692 703520
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 429212 142866 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 142860 429252 142866
rect 429200 142802 429252 142808
rect 433338 80472 433394 80481
rect 433338 80407 433394 80416
rect 415400 79552 415452 79558
rect 415400 79494 415452 79500
rect 397458 79112 397514 79121
rect 397458 79047 397514 79056
rect 192760 79008 192812 79014
rect 192760 78950 192812 78956
rect 233240 77172 233292 77178
rect 233240 77114 233292 77120
rect 222936 77104 222988 77110
rect 222936 77046 222988 77052
rect 220820 75744 220872 75750
rect 220820 75686 220872 75692
rect 195244 71664 195296 71670
rect 195244 71606 195296 71612
rect 195256 69018 195284 71606
rect 202328 70236 202380 70242
rect 202328 70178 202380 70184
rect 195244 69012 195296 69018
rect 195244 68954 195296 68960
rect 201132 69012 201184 69018
rect 201132 68954 201184 68960
rect 193220 68876 193272 68882
rect 193220 68818 193272 68824
rect 192576 60716 192628 60722
rect 192576 60658 192628 60664
rect 186332 16546 186912 16574
rect 187712 16546 188568 16574
rect 191852 16546 192064 16574
rect 184952 6886 185072 6914
rect 184952 480 184980 6886
rect 185584 3664 185636 3670
rect 185584 3606 185636 3612
rect 185596 3058 185624 3606
rect 186136 3324 186188 3330
rect 186136 3266 186188 3272
rect 185584 3052 185636 3058
rect 185584 2994 185636 3000
rect 186148 480 186176 3266
rect 182518 354 182630 480
rect 182192 326 182630 354
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188540 480 188568 16546
rect 190460 14272 190512 14278
rect 190460 14214 190512 14220
rect 189724 3392 189776 3398
rect 189724 3334 189776 3340
rect 189736 480 189764 3334
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 14214
rect 192036 480 192064 16546
rect 193232 480 193260 68818
rect 201144 66230 201172 68954
rect 201132 66224 201184 66230
rect 201132 66166 201184 66172
rect 202340 66162 202368 70178
rect 211068 69556 211120 69562
rect 211068 69498 211120 69504
rect 211080 67250 211108 69498
rect 211068 67244 211120 67250
rect 211068 67186 211120 67192
rect 203524 66224 203576 66230
rect 203524 66166 203576 66172
rect 202328 66156 202380 66162
rect 202328 66098 202380 66104
rect 200118 63064 200174 63073
rect 200118 62999 200174 63008
rect 197360 62824 197412 62830
rect 197360 62766 197412 62772
rect 194600 32632 194652 32638
rect 194600 32574 194652 32580
rect 193312 26988 193364 26994
rect 193312 26930 193364 26936
rect 193324 16574 193352 26930
rect 194612 16574 194640 32574
rect 197372 16574 197400 62766
rect 198740 32564 198792 32570
rect 198740 32506 198792 32512
rect 193324 16546 194456 16574
rect 194612 16546 195192 16574
rect 197372 16546 197952 16574
rect 194428 480 194456 16546
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 196808 6112 196860 6118
rect 196808 6054 196860 6060
rect 196820 480 196848 6054
rect 197924 480 197952 16546
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 32506
rect 200132 16574 200160 62999
rect 203536 55894 203564 66166
rect 205364 66156 205416 66162
rect 205364 66098 205416 66104
rect 205376 59362 205404 66098
rect 205364 59356 205416 59362
rect 205364 59298 205416 59304
rect 210424 59356 210476 59362
rect 210424 59298 210476 59304
rect 203524 55888 203576 55894
rect 203524 55830 203576 55836
rect 210436 51678 210464 59298
rect 210424 51672 210476 51678
rect 210424 51614 210476 51620
rect 212540 51672 212592 51678
rect 212540 51614 212592 51620
rect 209780 28212 209832 28218
rect 209780 28154 209832 28160
rect 205640 28144 205692 28150
rect 205640 28086 205692 28092
rect 201500 28076 201552 28082
rect 201500 28018 201552 28024
rect 200132 16546 200344 16574
rect 200316 480 200344 16546
rect 201512 11694 201540 28018
rect 201590 25528 201646 25537
rect 201590 25463 201646 25472
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 25463
rect 204260 23452 204312 23458
rect 204260 23394 204312 23400
rect 204272 16574 204300 23394
rect 205652 16574 205680 28086
rect 208400 23384 208452 23390
rect 208400 23326 208452 23332
rect 208412 16574 208440 23326
rect 204272 16546 205128 16574
rect 205652 16546 206232 16574
rect 208412 16546 208624 16574
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 203892 6860 203944 6866
rect 203892 6802 203944 6808
rect 203904 480 203932 6802
rect 205100 480 205128 16546
rect 206204 480 206232 16546
rect 207388 9240 207440 9246
rect 207388 9182 207440 9188
rect 207400 480 207428 9182
rect 208596 480 208624 16546
rect 209792 480 209820 28154
rect 211160 23316 211212 23322
rect 211160 23258 211212 23264
rect 211172 16574 211200 23258
rect 212552 16574 212580 51614
rect 216678 34232 216734 34241
rect 216678 34167 216734 34176
rect 215298 23352 215354 23361
rect 215298 23287 215354 23296
rect 211172 16546 211752 16574
rect 212552 16546 213408 16574
rect 210976 9172 211028 9178
rect 210976 9114 211028 9120
rect 210988 480 211016 9114
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213380 480 213408 16546
rect 214472 12436 214524 12442
rect 214472 12378 214524 12384
rect 214484 480 214512 12378
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 23287
rect 216692 16574 216720 34167
rect 218060 18692 218112 18698
rect 218060 18634 218112 18640
rect 216692 16546 216904 16574
rect 216876 480 216904 16546
rect 218072 3398 218100 18634
rect 220832 16574 220860 75686
rect 222948 68950 222976 77046
rect 230480 74520 230532 74526
rect 230480 74462 230532 74468
rect 226524 73772 226576 73778
rect 226524 73714 226576 73720
rect 226432 73704 226484 73710
rect 226432 73646 226484 73652
rect 226340 70304 226392 70310
rect 226340 70246 226392 70252
rect 224960 69624 225012 69630
rect 224960 69566 225012 69572
rect 222936 68944 222988 68950
rect 222936 68886 222988 68892
rect 224972 66978 225000 69566
rect 226352 67318 226380 70246
rect 226444 70242 226472 73646
rect 226432 70236 226484 70242
rect 226432 70178 226484 70184
rect 226536 69630 226564 73714
rect 226524 69624 226576 69630
rect 226524 69566 226576 69572
rect 226340 67312 226392 67318
rect 226340 67254 226392 67260
rect 224960 66972 225012 66978
rect 224960 66914 225012 66920
rect 223580 60240 223632 60246
rect 223580 60182 223632 60188
rect 220832 16546 221136 16574
rect 218150 6080 218206 6089
rect 218150 6015 218206 6024
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 218164 3074 218192 6015
rect 220452 5024 220504 5030
rect 220452 4966 220504 4972
rect 219256 3392 219308 3398
rect 219256 3334 219308 3340
rect 218072 3046 218192 3074
rect 218072 480 218100 3046
rect 219268 480 219296 3334
rect 220464 480 220492 4966
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 354 221136 16546
rect 222752 12368 222804 12374
rect 222752 12310 222804 12316
rect 222764 480 222792 12310
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 60182
rect 228364 55888 228416 55894
rect 228364 55830 228416 55836
rect 228376 44946 228404 55830
rect 228364 44940 228416 44946
rect 228364 44882 228416 44888
rect 226340 17672 226392 17678
rect 226340 17614 226392 17620
rect 226352 11694 226380 17614
rect 230492 16574 230520 74462
rect 230848 70372 230900 70378
rect 230848 70314 230900 70320
rect 230860 67182 230888 70314
rect 230848 67176 230900 67182
rect 230848 67118 230900 67124
rect 233252 16574 233280 77114
rect 303618 77072 303674 77081
rect 259460 77036 259512 77042
rect 303618 77007 303674 77016
rect 259460 76978 259512 76984
rect 256700 75676 256752 75682
rect 256700 75618 256752 75624
rect 242808 74452 242860 74458
rect 242808 74394 242860 74400
rect 242820 68882 242848 74394
rect 248972 74384 249024 74390
rect 248972 74326 249024 74332
rect 244372 74316 244424 74322
rect 244372 74258 244424 74264
rect 244280 72276 244332 72282
rect 244280 72218 244332 72224
rect 244292 69902 244320 72218
rect 244280 69896 244332 69902
rect 244280 69838 244332 69844
rect 242808 68876 242860 68882
rect 242808 68818 242860 68824
rect 244384 64874 244412 74258
rect 248984 67386 249012 74326
rect 251178 74080 251234 74089
rect 251178 74015 251234 74024
rect 248972 67380 249024 67386
rect 248972 67322 249024 67328
rect 244292 64846 244412 64874
rect 233884 44940 233936 44946
rect 233884 44882 233936 44888
rect 233896 40730 233924 44882
rect 233884 40724 233936 40730
rect 233884 40666 233936 40672
rect 241518 20496 241574 20505
rect 241518 20431 241574 20440
rect 237380 19916 237432 19922
rect 237380 19858 237432 19864
rect 234618 18592 234674 18601
rect 234618 18527 234674 18536
rect 230492 16546 231072 16574
rect 233252 16546 233464 16574
rect 226432 12300 226484 12306
rect 226432 12242 226484 12248
rect 226340 11688 226392 11694
rect 226340 11630 226392 11636
rect 226444 6914 226472 12242
rect 229376 12232 229428 12238
rect 229376 12174 229428 12180
rect 227536 11688 227588 11694
rect 227536 11630 227588 11636
rect 226352 6886 226472 6914
rect 225144 4140 225196 4146
rect 225144 4082 225196 4088
rect 225156 480 225184 4082
rect 226352 480 226380 6886
rect 227548 480 227576 11630
rect 228732 4072 228784 4078
rect 228732 4014 228784 4020
rect 228744 480 228772 4014
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229388 354 229416 12174
rect 231044 480 231072 16546
rect 232226 4040 232282 4049
rect 232226 3975 232282 3984
rect 232240 480 232268 3975
rect 233436 480 233464 16546
rect 234632 480 234660 18527
rect 237392 16574 237420 19858
rect 241532 16574 241560 20431
rect 244292 16574 244320 64846
rect 245660 40724 245712 40730
rect 245660 40666 245712 40672
rect 245672 36650 245700 40666
rect 245660 36644 245712 36650
rect 245660 36586 245712 36592
rect 237392 16546 237696 16574
rect 241532 16546 241744 16574
rect 244292 16546 245240 16574
rect 236550 10432 236606 10441
rect 236550 10367 236606 10376
rect 235814 3904 235870 3913
rect 235814 3839 235870 3848
rect 235828 480 235856 3839
rect 229806 354 229918 480
rect 229388 326 229918 354
rect 229806 -960 229918 326
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 10367
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 240140 12164 240192 12170
rect 240140 12106 240192 12112
rect 239312 4004 239364 4010
rect 239312 3946 239364 3952
rect 239324 480 239352 3946
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 12106
rect 241716 480 241744 16546
rect 242900 12096 242952 12102
rect 242900 12038 242952 12044
rect 242912 3398 242940 12038
rect 242990 3768 243046 3777
rect 242990 3703 243046 3712
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 243004 1850 243032 3703
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 242912 1822 243032 1850
rect 242912 480 242940 1822
rect 244108 480 244136 3334
rect 245212 480 245240 16546
rect 248420 15972 248472 15978
rect 248420 15914 248472 15920
rect 247592 9104 247644 9110
rect 247592 9046 247644 9052
rect 246396 6792 246448 6798
rect 246396 6734 246448 6740
rect 246408 480 246436 6734
rect 247604 480 247632 9046
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 15914
rect 249982 6896 250038 6905
rect 249982 6831 250038 6840
rect 249996 480 250024 6831
rect 251192 4010 251220 74015
rect 255320 73092 255372 73098
rect 255320 73034 255372 73040
rect 255332 71670 255360 73034
rect 255320 71664 255372 71670
rect 255320 71606 255372 71612
rect 254584 70168 254636 70174
rect 254584 70110 254636 70116
rect 254596 64054 254624 70110
rect 254584 64048 254636 64054
rect 254584 63990 254636 63996
rect 253940 26036 253992 26042
rect 253940 25978 253992 25984
rect 253952 16574 253980 25978
rect 255320 20664 255372 20670
rect 255320 20606 255372 20612
rect 255332 16574 255360 20606
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 251270 12064 251326 12073
rect 251270 11999 251326 12008
rect 251180 4004 251232 4010
rect 251180 3946 251232 3952
rect 251284 3482 251312 11999
rect 253478 6760 253534 6769
rect 253478 6695 253534 6704
rect 252376 4004 252428 4010
rect 252376 3946 252428 3952
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3946
rect 253492 480 253520 6695
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 256712 354 256740 75618
rect 256792 74248 256844 74254
rect 256792 74190 256844 74196
rect 256804 70174 256832 74190
rect 257344 71596 257396 71602
rect 257344 71538 257396 71544
rect 256792 70168 256844 70174
rect 256792 70110 256844 70116
rect 257356 60246 257384 71538
rect 257344 60240 257396 60246
rect 257344 60182 257396 60188
rect 259472 11694 259500 76978
rect 273536 76968 273588 76974
rect 273536 76910 273588 76916
rect 267740 76900 267792 76906
rect 267740 76842 267792 76848
rect 262864 75608 262916 75614
rect 262864 75550 262916 75556
rect 261484 74180 261536 74186
rect 261484 74122 261536 74128
rect 260196 71528 260248 71534
rect 260196 71470 260248 71476
rect 259552 67380 259604 67386
rect 259552 67322 259604 67328
rect 259564 63578 259592 67322
rect 260208 66230 260236 71470
rect 260196 66224 260248 66230
rect 260196 66166 260248 66172
rect 260472 64048 260524 64054
rect 260472 63990 260524 63996
rect 259552 63572 259604 63578
rect 259552 63514 259604 63520
rect 260484 59362 260512 63990
rect 261496 62898 261524 74122
rect 261574 71768 261630 71777
rect 261574 71703 261630 71712
rect 261484 62892 261536 62898
rect 261484 62834 261536 62840
rect 261588 62830 261616 71703
rect 262876 67590 262904 75550
rect 264980 72412 265032 72418
rect 264980 72354 265032 72360
rect 263048 70100 263100 70106
rect 263048 70042 263100 70048
rect 262864 67584 262916 67590
rect 262864 67526 262916 67532
rect 263060 63782 263088 70042
rect 264992 67386 265020 72354
rect 265624 70032 265676 70038
rect 265624 69974 265676 69980
rect 264980 67380 265032 67386
rect 264980 67322 265032 67328
rect 263508 66224 263560 66230
rect 263508 66166 263560 66172
rect 263048 63776 263100 63782
rect 263048 63718 263100 63724
rect 263416 63572 263468 63578
rect 263416 63514 263468 63520
rect 261576 62824 261628 62830
rect 261576 62766 261628 62772
rect 261484 60240 261536 60246
rect 261484 60182 261536 60188
rect 260472 59356 260524 59362
rect 260472 59298 260524 59304
rect 261496 53106 261524 60182
rect 262220 59356 262272 59362
rect 262220 59298 262272 59304
rect 262232 56574 262260 59298
rect 263428 57254 263456 63514
rect 263520 59362 263548 66166
rect 265440 63776 265492 63782
rect 265440 63718 265492 63724
rect 265452 60654 265480 63718
rect 265440 60648 265492 60654
rect 265440 60590 265492 60596
rect 263508 59356 263560 59362
rect 263508 59298 263560 59304
rect 263416 57248 263468 57254
rect 263416 57190 263468 57196
rect 262220 56568 262272 56574
rect 262220 56510 262272 56516
rect 265636 53174 265664 69974
rect 267004 67584 267056 67590
rect 267004 67526 267056 67532
rect 266360 56568 266412 56574
rect 266360 56510 266412 56516
rect 266372 53242 266400 56510
rect 267016 54534 267044 67526
rect 267004 54528 267056 54534
rect 267004 54470 267056 54476
rect 266360 53236 266412 53242
rect 266360 53178 266412 53184
rect 265624 53168 265676 53174
rect 265624 53110 265676 53116
rect 261484 53100 261536 53106
rect 261484 53042 261536 53048
rect 259552 20596 259604 20602
rect 259552 20538 259604 20544
rect 259460 11688 259512 11694
rect 259460 11630 259512 11636
rect 259564 6914 259592 20538
rect 262220 20528 262272 20534
rect 262220 20470 262272 20476
rect 262232 16574 262260 20470
rect 266358 20360 266414 20369
rect 266358 20295 266414 20304
rect 266372 16574 266400 20295
rect 267752 16574 267780 76842
rect 272890 75712 272946 75721
rect 272890 75647 272946 75656
rect 272904 71466 272932 75647
rect 273548 71806 273576 76910
rect 280344 76832 280396 76838
rect 280344 76774 280396 76780
rect 280356 75818 280384 76774
rect 280344 75812 280396 75818
rect 280344 75754 280396 75760
rect 283196 75812 283248 75818
rect 283196 75754 283248 75760
rect 274640 75540 274692 75546
rect 274640 75482 274692 75488
rect 273536 71800 273588 71806
rect 273536 71742 273588 71748
rect 272524 71460 272576 71466
rect 272524 71402 272576 71408
rect 272892 71460 272944 71466
rect 272892 71402 272944 71408
rect 271144 69964 271196 69970
rect 271144 69906 271196 69912
rect 269856 68808 269908 68814
rect 269856 68750 269908 68756
rect 269120 67244 269172 67250
rect 269120 67186 269172 67192
rect 269132 63918 269160 67186
rect 269120 63912 269172 63918
rect 269120 63854 269172 63860
rect 269868 60654 269896 68750
rect 269764 60648 269816 60654
rect 269764 60590 269816 60596
rect 269856 60648 269908 60654
rect 269856 60590 269908 60596
rect 268844 59356 268896 59362
rect 268844 59298 268896 59304
rect 268856 56574 268884 59298
rect 268844 56568 268896 56574
rect 268844 56510 268896 56516
rect 269776 47598 269804 60590
rect 271156 55894 271184 69906
rect 271604 67040 271656 67046
rect 271604 66982 271656 66988
rect 271616 62082 271644 66982
rect 271880 63912 271932 63918
rect 271880 63854 271932 63860
rect 271604 62076 271656 62082
rect 271604 62018 271656 62024
rect 271892 58886 271920 63854
rect 272536 58954 272564 71402
rect 273996 70236 274048 70242
rect 273996 70178 274048 70184
rect 273444 67380 273496 67386
rect 273444 67322 273496 67328
rect 272524 58948 272576 58954
rect 272524 58890 272576 58896
rect 271880 58880 271932 58886
rect 271880 58822 271932 58828
rect 273456 58818 273484 67322
rect 273444 58812 273496 58818
rect 273444 58754 273496 58760
rect 273260 57248 273312 57254
rect 273260 57190 273312 57196
rect 271144 55888 271196 55894
rect 271144 55830 271196 55836
rect 273272 54602 273300 57190
rect 273260 54596 273312 54602
rect 273260 54538 273312 54544
rect 272524 53168 272576 53174
rect 272524 53110 272576 53116
rect 269764 47592 269816 47598
rect 269764 47534 269816 47540
rect 272536 23322 272564 53110
rect 273904 53100 273956 53106
rect 273904 53042 273956 53048
rect 273916 36718 273944 53042
rect 274008 53038 274036 70178
rect 274088 69624 274140 69630
rect 274088 69566 274140 69572
rect 274100 53174 274128 69566
rect 274272 56568 274324 56574
rect 274272 56510 274324 56516
rect 274088 53168 274140 53174
rect 274088 53110 274140 53116
rect 273996 53032 274048 53038
rect 273996 52974 274048 52980
rect 274284 52970 274312 56510
rect 274272 52964 274324 52970
rect 274272 52906 274324 52912
rect 273904 36712 273956 36718
rect 273904 36654 273956 36660
rect 273996 36644 274048 36650
rect 273996 36586 274048 36592
rect 274008 24206 274036 36586
rect 273996 24200 274048 24206
rect 273996 24142 274048 24148
rect 272524 23316 272576 23322
rect 272524 23258 272576 23264
rect 273260 23248 273312 23254
rect 273260 23190 273312 23196
rect 269120 20460 269172 20466
rect 269120 20402 269172 20408
rect 269132 16574 269160 20402
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 267752 16546 268424 16574
rect 269132 16546 270080 16574
rect 261760 14340 261812 14346
rect 261760 14282 261812 14288
rect 260656 11688 260708 11694
rect 260656 11630 260708 11636
rect 259472 6886 259592 6914
rect 258264 3936 258316 3942
rect 258264 3878 258316 3884
rect 258276 480 258304 3878
rect 259472 480 259500 6886
rect 260668 480 260696 11630
rect 261772 480 261800 14282
rect 257038 354 257150 480
rect 256712 326 257150 354
rect 257038 -960 257150 326
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264980 14408 265032 14414
rect 264980 14350 265032 14356
rect 264150 3632 264206 3641
rect 264150 3567 264206 3576
rect 264164 480 264192 3567
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 14350
rect 266556 480 266584 16546
rect 267740 6724 267792 6730
rect 267740 6666 267792 6672
rect 267752 480 267780 6666
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 272430 11928 272486 11937
rect 272430 11863 272486 11872
rect 271234 6624 271290 6633
rect 271234 6559 271290 6568
rect 271248 480 271276 6559
rect 272444 480 272472 11863
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 23190
rect 274652 16574 274680 75482
rect 282184 74112 282236 74118
rect 282184 74054 282236 74060
rect 281816 74044 281868 74050
rect 281816 73986 281868 73992
rect 281356 73024 281408 73030
rect 281356 72966 281408 72972
rect 275284 72344 275336 72350
rect 275284 72286 275336 72292
rect 274732 60648 274784 60654
rect 274732 60590 274784 60596
rect 274744 56982 274772 60590
rect 274732 56976 274784 56982
rect 274732 56918 274784 56924
rect 275296 50386 275324 72286
rect 276020 71800 276072 71806
rect 276020 71742 276072 71748
rect 276032 67046 276060 71742
rect 280894 71632 280950 71641
rect 280894 71567 280950 71576
rect 280804 70168 280856 70174
rect 280804 70110 280856 70116
rect 279424 67312 279476 67318
rect 279424 67254 279476 67260
rect 276020 67040 276072 67046
rect 276020 66982 276072 66988
rect 276664 62892 276716 62898
rect 276664 62834 276716 62840
rect 276112 54596 276164 54602
rect 276112 54538 276164 54544
rect 276020 52964 276072 52970
rect 276020 52906 276072 52912
rect 276032 50454 276060 52906
rect 276020 50448 276072 50454
rect 276020 50390 276072 50396
rect 275284 50380 275336 50386
rect 275284 50322 275336 50328
rect 276124 47666 276152 54538
rect 276676 47734 276704 62834
rect 277952 62076 278004 62082
rect 277952 62018 278004 62024
rect 277964 58614 277992 62018
rect 277952 58608 278004 58614
rect 277952 58550 278004 58556
rect 279436 57254 279464 67254
rect 280816 62082 280844 70110
rect 280908 62898 280936 71567
rect 280988 71392 281040 71398
rect 280988 71334 281040 71340
rect 281000 62966 281028 71334
rect 281368 69970 281396 72966
rect 281448 72956 281500 72962
rect 281448 72898 281500 72904
rect 281356 69964 281408 69970
rect 281356 69906 281408 69912
rect 281460 69018 281488 72898
rect 281448 69012 281500 69018
rect 281448 68954 281500 68960
rect 281828 68814 281856 73986
rect 282000 72888 282052 72894
rect 282000 72830 282052 72836
rect 281908 72820 281960 72826
rect 281908 72762 281960 72768
rect 281920 69290 281948 72762
rect 281908 69284 281960 69290
rect 281908 69226 281960 69232
rect 282012 69222 282040 72830
rect 282000 69216 282052 69222
rect 282000 69158 282052 69164
rect 281816 68808 281868 68814
rect 281816 68750 281868 68756
rect 282196 63510 282224 74054
rect 283208 71738 283236 75754
rect 290464 73976 290516 73982
rect 290464 73918 290516 73924
rect 295338 73944 295394 73953
rect 289174 72584 289230 72593
rect 289174 72519 289230 72528
rect 283196 71732 283248 71738
rect 283196 71674 283248 71680
rect 284300 71460 284352 71466
rect 284300 71402 284352 71408
rect 284312 67046 284340 71402
rect 285772 69964 285824 69970
rect 285772 69906 285824 69912
rect 284392 69284 284444 69290
rect 284392 69226 284444 69232
rect 282276 67040 282328 67046
rect 282276 66982 282328 66988
rect 284300 67040 284352 67046
rect 284300 66982 284352 66988
rect 282288 64122 282316 66982
rect 284404 65686 284432 69226
rect 284484 69216 284536 69222
rect 284484 69158 284536 69164
rect 284392 65680 284444 65686
rect 284392 65622 284444 65628
rect 284496 65618 284524 69158
rect 285680 67108 285732 67114
rect 285680 67050 285732 67056
rect 284484 65612 284536 65618
rect 284484 65554 284536 65560
rect 285692 64326 285720 67050
rect 285784 64938 285812 69906
rect 285772 64932 285824 64938
rect 285772 64874 285824 64880
rect 289084 64932 289136 64938
rect 289084 64874 289136 64880
rect 285680 64320 285732 64326
rect 285680 64262 285732 64268
rect 282276 64116 282328 64122
rect 282276 64058 282328 64064
rect 282184 63504 282236 63510
rect 282184 63446 282236 63452
rect 287888 63504 287940 63510
rect 287888 63446 287940 63452
rect 280988 62960 281040 62966
rect 280988 62902 281040 62908
rect 280896 62892 280948 62898
rect 280896 62834 280948 62840
rect 284300 62824 284352 62830
rect 284300 62766 284352 62772
rect 280804 62076 280856 62082
rect 280804 62018 280856 62024
rect 280988 58948 281040 58954
rect 280988 58890 281040 58896
rect 279424 57248 279476 57254
rect 279424 57190 279476 57196
rect 277768 56976 277820 56982
rect 277768 56918 277820 56924
rect 277780 49706 277808 56918
rect 281000 56574 281028 58890
rect 284312 58818 284340 62766
rect 287704 62076 287756 62082
rect 287704 62018 287756 62024
rect 286416 58880 286468 58886
rect 286416 58822 286468 58828
rect 283748 58812 283800 58818
rect 283748 58754 283800 58760
rect 284300 58812 284352 58818
rect 284300 58754 284352 58760
rect 283564 58608 283616 58614
rect 283564 58550 283616 58556
rect 280988 56568 281040 56574
rect 280988 56510 281040 56516
rect 280804 53236 280856 53242
rect 280804 53178 280856 53184
rect 277768 49700 277820 49706
rect 277768 49642 277820 49648
rect 276664 47728 276716 47734
rect 276664 47670 276716 47676
rect 276112 47660 276164 47666
rect 276112 47602 276164 47608
rect 280816 26042 280844 53178
rect 282920 49700 282972 49706
rect 282920 49642 282972 49648
rect 282184 47728 282236 47734
rect 282184 47670 282236 47676
rect 280804 26036 280856 26042
rect 280804 25978 280856 25984
rect 275008 23316 275060 23322
rect 275008 23258 275060 23264
rect 275020 20466 275048 23258
rect 280160 23180 280212 23186
rect 280160 23122 280212 23128
rect 275008 20460 275060 20466
rect 275008 20402 275060 20408
rect 276020 20392 276072 20398
rect 276020 20334 276072 20340
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 3942 276060 20334
rect 280172 16574 280200 23122
rect 280172 16546 280752 16574
rect 276112 15156 276164 15162
rect 276112 15098 276164 15104
rect 276020 3936 276072 3942
rect 276020 3878 276072 3884
rect 276124 3482 276152 15098
rect 279056 15088 279108 15094
rect 279056 15030 279108 15036
rect 278320 6656 278372 6662
rect 278320 6598 278372 6604
rect 276756 3936 276808 3942
rect 276756 3878 276808 3884
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 3878
rect 278332 480 278360 6598
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 15030
rect 280724 480 280752 16546
rect 282196 9110 282224 47670
rect 282932 46238 282960 49642
rect 282920 46232 282972 46238
rect 282920 46174 282972 46180
rect 283576 26178 283604 58550
rect 283656 47592 283708 47598
rect 283656 47534 283708 47540
rect 283564 26172 283616 26178
rect 283564 26114 283616 26120
rect 283668 26110 283696 47534
rect 283760 36786 283788 58754
rect 286324 56568 286376 56574
rect 286324 56510 286376 56516
rect 284300 54528 284352 54534
rect 284300 54470 284352 54476
rect 284312 51746 284340 54470
rect 284300 51740 284352 51746
rect 284300 51682 284352 51688
rect 285680 50380 285732 50386
rect 285680 50322 285732 50328
rect 284944 47660 284996 47666
rect 284944 47602 284996 47608
rect 284956 45558 284984 47602
rect 285692 47598 285720 50322
rect 285680 47592 285732 47598
rect 285680 47534 285732 47540
rect 284944 45552 284996 45558
rect 284944 45494 284996 45500
rect 286336 44470 286364 56510
rect 286428 49162 286456 58822
rect 287060 57248 287112 57254
rect 287060 57190 287112 57196
rect 287072 54534 287100 57190
rect 287060 54528 287112 54534
rect 287060 54470 287112 54476
rect 287716 54126 287744 62018
rect 287900 59702 287928 63446
rect 287888 59696 287940 59702
rect 287888 59638 287940 59644
rect 287704 54120 287756 54126
rect 287704 54062 287756 54068
rect 287612 50448 287664 50454
rect 287612 50390 287664 50396
rect 286416 49156 286468 49162
rect 286416 49098 286468 49104
rect 287624 48278 287652 50390
rect 287612 48272 287664 48278
rect 287612 48214 287664 48220
rect 287612 45552 287664 45558
rect 287612 45494 287664 45500
rect 286324 44464 286376 44470
rect 286324 44406 286376 44412
rect 287624 42430 287652 45494
rect 287612 42424 287664 42430
rect 287612 42366 287664 42372
rect 289096 42158 289124 64874
rect 289188 60382 289216 72519
rect 289360 71732 289412 71738
rect 289360 71674 289412 71680
rect 289372 68270 289400 71674
rect 289360 68264 289412 68270
rect 289360 68206 289412 68212
rect 289360 64116 289412 64122
rect 289360 64058 289412 64064
rect 289372 60858 289400 64058
rect 289360 60852 289412 60858
rect 289360 60794 289412 60800
rect 289176 60376 289228 60382
rect 289176 60318 289228 60324
rect 290476 50590 290504 73918
rect 295338 73879 295394 73888
rect 295984 73908 296036 73914
rect 295352 72826 295380 73879
rect 295984 73850 296036 73856
rect 295340 72820 295392 72826
rect 295340 72762 295392 72768
rect 294604 68944 294656 68950
rect 294604 68886 294656 68892
rect 294616 64394 294644 68886
rect 294604 64388 294656 64394
rect 294604 64330 294656 64336
rect 294052 64320 294104 64326
rect 294052 64262 294104 64268
rect 291936 60852 291988 60858
rect 291936 60794 291988 60800
rect 290556 59696 290608 59702
rect 290556 59638 290608 59644
rect 290464 50584 290516 50590
rect 290464 50526 290516 50532
rect 290568 50386 290596 59638
rect 291844 55888 291896 55894
rect 291844 55830 291896 55836
rect 290832 51740 290884 51746
rect 290832 51682 290884 51688
rect 290556 50380 290608 50386
rect 290556 50322 290608 50328
rect 290844 49094 290872 51682
rect 290832 49088 290884 49094
rect 290832 49030 290884 49036
rect 290648 46232 290700 46238
rect 290648 46174 290700 46180
rect 289728 44464 289780 44470
rect 289728 44406 289780 44412
rect 289084 42152 289136 42158
rect 289084 42094 289136 42100
rect 283748 36780 283800 36786
rect 283748 36722 283800 36728
rect 284944 36712 284996 36718
rect 284944 36654 284996 36660
rect 283656 26104 283708 26110
rect 283656 26046 283708 26052
rect 284956 24138 284984 36654
rect 289740 36650 289768 44406
rect 290660 40050 290688 46174
rect 290648 40044 290700 40050
rect 290648 39986 290700 39992
rect 290372 36780 290424 36786
rect 290372 36722 290424 36728
rect 289728 36644 289780 36650
rect 289728 36586 289780 36592
rect 290384 29714 290412 36722
rect 290372 29708 290424 29714
rect 290372 29650 290424 29656
rect 289820 28960 289872 28966
rect 289820 28902 289872 28908
rect 284944 24132 284996 24138
rect 284944 24074 284996 24080
rect 284298 23216 284354 23225
rect 284298 23151 284354 23160
rect 283104 15020 283156 15026
rect 283104 14962 283156 14968
rect 282184 9104 282236 9110
rect 282184 9046 282236 9052
rect 281908 6588 281960 6594
rect 281908 6530 281960 6536
rect 281920 480 281948 6530
rect 283116 480 283144 14962
rect 284312 480 284340 23151
rect 287058 23080 287114 23089
rect 287058 23015 287114 23024
rect 287072 16574 287100 23015
rect 288348 20460 288400 20466
rect 288348 20402 288400 20408
rect 288360 17746 288388 20402
rect 288348 17740 288400 17746
rect 288348 17682 288400 17688
rect 287072 16546 287376 16574
rect 286598 14512 286654 14521
rect 286598 14447 286654 14456
rect 285402 6488 285458 6497
rect 285402 6423 285458 6432
rect 285416 480 285444 6423
rect 286612 480 286640 14447
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 288990 6352 289046 6361
rect 288990 6287 289046 6296
rect 289004 480 289032 6287
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 28902
rect 291856 24614 291884 55830
rect 291948 54194 291976 60794
rect 293960 60376 294012 60382
rect 293960 60318 294012 60324
rect 293972 55894 294000 60318
rect 294064 60246 294092 64262
rect 294052 60240 294104 60246
rect 294052 60182 294104 60188
rect 293960 55888 294012 55894
rect 293960 55830 294012 55836
rect 291936 54188 291988 54194
rect 291936 54130 291988 54136
rect 295340 54120 295392 54126
rect 295340 54062 295392 54068
rect 293224 50584 293276 50590
rect 293224 50526 293276 50532
rect 291936 48272 291988 48278
rect 291936 48214 291988 48220
rect 291844 24608 291896 24614
rect 291844 24550 291896 24556
rect 291200 23112 291252 23118
rect 291200 23054 291252 23060
rect 291212 16574 291240 23054
rect 291948 22914 291976 48214
rect 292028 42424 292080 42430
rect 292028 42366 292080 42372
rect 292040 24274 292068 42366
rect 293236 42090 293264 50526
rect 295352 49298 295380 54062
rect 295996 53242 296024 73850
rect 300308 72820 300360 72826
rect 300308 72762 300360 72768
rect 299388 72752 299440 72758
rect 299388 72694 299440 72700
rect 297364 71664 297416 71670
rect 297364 71606 297416 71612
rect 297376 62150 297404 71606
rect 299400 69970 299428 72694
rect 299388 69964 299440 69970
rect 299388 69906 299440 69912
rect 298744 69012 298796 69018
rect 298744 68954 298796 68960
rect 297364 62144 297416 62150
rect 297364 62086 297416 62092
rect 295984 53236 296036 53242
rect 295984 53178 296036 53184
rect 297364 53168 297416 53174
rect 297364 53110 297416 53116
rect 295340 49292 295392 49298
rect 295340 49234 295392 49240
rect 294604 49156 294656 49162
rect 294604 49098 294656 49104
rect 293868 47592 293920 47598
rect 293868 47534 293920 47540
rect 293880 45014 293908 47534
rect 293868 45008 293920 45014
rect 293868 44950 293920 44956
rect 294616 44946 294644 49098
rect 294604 44940 294656 44946
rect 294604 44882 294656 44888
rect 297376 42838 297404 53110
rect 297456 53100 297508 53106
rect 297456 53042 297508 53048
rect 297468 42906 297496 53042
rect 298756 44742 298784 68954
rect 300124 65680 300176 65686
rect 300124 65622 300176 65628
rect 299112 54188 299164 54194
rect 299112 54130 299164 54136
rect 299124 49842 299152 54130
rect 299112 49836 299164 49842
rect 299112 49778 299164 49784
rect 300136 49162 300164 65622
rect 300216 65612 300268 65618
rect 300216 65554 300268 65560
rect 300228 49230 300256 65554
rect 300320 56574 300348 72762
rect 300400 68740 300452 68746
rect 300400 68682 300452 68688
rect 300412 63170 300440 68682
rect 303160 68672 303212 68678
rect 303160 68614 303212 68620
rect 300492 68264 300544 68270
rect 300492 68206 300544 68212
rect 300400 63164 300452 63170
rect 300400 63106 300452 63112
rect 300504 63102 300532 68206
rect 302976 67040 303028 67046
rect 302976 66982 303028 66988
rect 301504 64388 301556 64394
rect 301504 64330 301556 64336
rect 300492 63096 300544 63102
rect 300492 63038 300544 63044
rect 301516 61402 301544 64330
rect 302332 62960 302384 62966
rect 302332 62902 302384 62908
rect 302240 62892 302292 62898
rect 302240 62834 302292 62840
rect 301504 61396 301556 61402
rect 301504 61338 301556 61344
rect 302252 59770 302280 62834
rect 302240 59764 302292 59770
rect 302240 59706 302292 59712
rect 302344 59634 302372 62902
rect 302884 62144 302936 62150
rect 302884 62086 302936 62092
rect 302332 59628 302384 59634
rect 302332 59570 302384 59576
rect 301320 58812 301372 58818
rect 301320 58754 301372 58760
rect 300308 56568 300360 56574
rect 300308 56510 300360 56516
rect 301332 56506 301360 58754
rect 302240 56568 302292 56574
rect 302240 56510 302292 56516
rect 301320 56500 301372 56506
rect 301320 56442 301372 56448
rect 302252 52018 302280 56510
rect 302240 52012 302292 52018
rect 302240 51954 302292 51960
rect 301504 49836 301556 49842
rect 301504 49778 301556 49784
rect 300216 49224 300268 49230
rect 300216 49166 300268 49172
rect 300124 49156 300176 49162
rect 300124 49098 300176 49104
rect 298744 44736 298796 44742
rect 298744 44678 298796 44684
rect 297456 42900 297508 42906
rect 297456 42842 297508 42848
rect 300768 42900 300820 42906
rect 300768 42842 300820 42848
rect 297364 42832 297416 42838
rect 297364 42774 297416 42780
rect 300124 42832 300176 42838
rect 300124 42774 300176 42780
rect 297640 42152 297692 42158
rect 297640 42094 297692 42100
rect 293224 42084 293276 42090
rect 293224 42026 293276 42032
rect 294604 40044 294656 40050
rect 294604 39986 294656 39992
rect 292578 28520 292634 28529
rect 292578 28455 292634 28464
rect 292028 24268 292080 24274
rect 292028 24210 292080 24216
rect 291936 22908 291988 22914
rect 291936 22850 291988 22856
rect 292592 16574 292620 28455
rect 292764 26172 292816 26178
rect 292764 26114 292816 26120
rect 292672 24200 292724 24206
rect 292672 24142 292724 24148
rect 292684 20466 292712 24142
rect 292672 20460 292724 20466
rect 292672 20402 292724 20408
rect 292776 20398 292804 26114
rect 294052 26104 294104 26110
rect 294052 26046 294104 26052
rect 293960 23044 294012 23050
rect 293960 22986 294012 22992
rect 292764 20392 292816 20398
rect 292764 20334 292816 20340
rect 293972 16574 294000 22986
rect 294064 18766 294092 26046
rect 294144 26036 294196 26042
rect 294144 25978 294196 25984
rect 294052 18760 294104 18766
rect 294052 18702 294104 18708
rect 294156 17678 294184 25978
rect 294328 24608 294380 24614
rect 294328 24550 294380 24556
rect 294340 22098 294368 24550
rect 294616 23050 294644 39986
rect 297652 37262 297680 42094
rect 297640 37256 297692 37262
rect 297640 37198 297692 37204
rect 300136 26994 300164 42774
rect 300492 37256 300544 37262
rect 300492 37198 300544 37204
rect 300504 30326 300532 37198
rect 300780 36106 300808 42842
rect 301516 39438 301544 49778
rect 302240 45008 302292 45014
rect 302240 44950 302292 44956
rect 301504 39432 301556 39438
rect 301504 39374 301556 39380
rect 302252 36718 302280 44950
rect 302240 36712 302292 36718
rect 302240 36654 302292 36660
rect 300768 36100 300820 36106
rect 300768 36042 300820 36048
rect 300492 30320 300544 30326
rect 300492 30262 300544 30268
rect 302240 30320 302292 30326
rect 302240 30262 302292 30268
rect 300124 26988 300176 26994
rect 300124 26930 300176 26936
rect 302252 26382 302280 30262
rect 302240 26376 302292 26382
rect 302240 26318 302292 26324
rect 302896 24886 302924 62086
rect 302988 36786 303016 66982
rect 303068 60240 303120 60246
rect 303068 60182 303120 60188
rect 303080 46238 303108 60182
rect 303172 57254 303200 68614
rect 303250 68368 303306 68377
rect 303250 68303 303306 68312
rect 303264 59362 303292 68303
rect 303252 59356 303304 59362
rect 303252 59298 303304 59304
rect 303160 57248 303212 57254
rect 303160 57190 303212 57196
rect 303528 55888 303580 55894
rect 303528 55830 303580 55836
rect 303540 51746 303568 55830
rect 303528 51740 303580 51746
rect 303528 51682 303580 51688
rect 303068 46232 303120 46238
rect 303068 46174 303120 46180
rect 302976 36780 303028 36786
rect 302976 36722 303028 36728
rect 302884 24880 302936 24886
rect 302884 24822 302936 24828
rect 300676 24268 300728 24274
rect 300676 24210 300728 24216
rect 294604 23044 294656 23050
rect 294604 22986 294656 22992
rect 294328 22092 294380 22098
rect 294328 22034 294380 22040
rect 298008 22092 298060 22098
rect 298008 22034 298060 22040
rect 298020 18698 298048 22034
rect 300688 20670 300716 24210
rect 300860 22976 300912 22982
rect 300860 22918 300912 22924
rect 300676 20664 300728 20670
rect 300676 20606 300728 20612
rect 300124 20460 300176 20466
rect 300124 20402 300176 20408
rect 298100 20324 298152 20330
rect 298100 20266 298152 20272
rect 298008 18692 298060 18698
rect 298008 18634 298060 18640
rect 297364 17740 297416 17746
rect 297364 17682 297416 17688
rect 294144 17672 294196 17678
rect 294144 17614 294196 17620
rect 291212 16546 291424 16574
rect 292592 16546 293264 16574
rect 293972 16546 294920 16574
rect 291396 480 291424 16546
rect 292580 6520 292632 6526
rect 292580 6462 292632 6468
rect 292592 480 292620 6462
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 297272 14952 297324 14958
rect 297272 14894 297324 14900
rect 296076 6452 296128 6458
rect 296076 6394 296128 6400
rect 296088 480 296116 6394
rect 297284 480 297312 14894
rect 297376 8294 297404 17682
rect 297364 8288 297416 8294
rect 297364 8230 297416 8236
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 20266
rect 300136 15026 300164 20402
rect 300872 16574 300900 22918
rect 303632 16574 303660 77007
rect 311900 76764 311952 76770
rect 311900 76706 311952 76712
rect 305642 75576 305698 75585
rect 311912 75546 311940 76706
rect 336740 76696 336792 76702
rect 336740 76638 336792 76644
rect 305642 75511 305698 75520
rect 311900 75540 311952 75546
rect 303712 63096 303764 63102
rect 303712 63038 303764 63044
rect 303724 60246 303752 63038
rect 303712 60240 303764 60246
rect 303712 60182 303764 60188
rect 305656 54602 305684 75511
rect 311900 75482 311952 75488
rect 320548 75540 320600 75546
rect 320548 75482 320600 75488
rect 310242 75440 310298 75449
rect 310242 75375 310298 75384
rect 305736 71324 305788 71330
rect 305736 71266 305788 71272
rect 305748 54670 305776 71266
rect 310256 70106 310284 75375
rect 318154 73808 318210 73817
rect 318154 73743 318210 73752
rect 311164 72684 311216 72690
rect 311164 72626 311216 72632
rect 310426 71496 310482 71505
rect 310426 71431 310482 71440
rect 310244 70100 310296 70106
rect 310244 70042 310296 70048
rect 309784 69964 309836 69970
rect 309784 69906 309836 69912
rect 307668 63164 307720 63170
rect 307668 63106 307720 63112
rect 306012 59764 306064 59770
rect 306012 59706 306064 59712
rect 305828 59356 305880 59362
rect 305828 59298 305880 59304
rect 305736 54664 305788 54670
rect 305736 54606 305788 54612
rect 305644 54596 305696 54602
rect 305644 54538 305696 54544
rect 305000 52012 305052 52018
rect 305000 51954 305052 51960
rect 304264 49292 304316 49298
rect 304264 49234 304316 49240
rect 303804 44736 303856 44742
rect 303804 44678 303856 44684
rect 303712 42084 303764 42090
rect 303712 42026 303764 42032
rect 303724 40050 303752 42026
rect 303712 40044 303764 40050
rect 303712 39986 303764 39992
rect 303816 37942 303844 44678
rect 303804 37936 303856 37942
rect 303804 37878 303856 37884
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 300124 15020 300176 15026
rect 300124 14962 300176 14968
rect 299664 6384 299716 6390
rect 299664 6326 299716 6332
rect 299676 480 299704 6326
rect 300768 6316 300820 6322
rect 300768 6258 300820 6264
rect 300780 480 300808 6258
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303158 9208 303214 9217
rect 303158 9143 303214 9152
rect 302148 9104 302200 9110
rect 302148 9046 302200 9052
rect 302160 3398 302188 9046
rect 302148 3392 302200 3398
rect 302148 3334 302200 3340
rect 303172 480 303200 9143
rect 303528 8288 303580 8294
rect 303528 8230 303580 8236
rect 303540 4078 303568 8230
rect 303528 4072 303580 4078
rect 303528 4014 303580 4020
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 304276 14958 304304 49234
rect 305012 47598 305040 51954
rect 305840 50454 305868 59298
rect 305920 56500 305972 56506
rect 305920 56442 305972 56448
rect 305828 50448 305880 50454
rect 305828 50390 305880 50396
rect 305932 50386 305960 56442
rect 306024 54738 306052 59706
rect 306104 59628 306156 59634
rect 306104 59570 306156 59576
rect 306116 54806 306144 59570
rect 307680 55894 307708 63106
rect 309796 56574 309824 69906
rect 310440 69562 310468 71431
rect 310428 69556 310480 69562
rect 310428 69498 310480 69504
rect 311176 61946 311204 72626
rect 318168 71330 318196 73743
rect 318156 71324 318208 71330
rect 318156 71266 318208 71272
rect 312544 70100 312596 70106
rect 312544 70042 312596 70048
rect 311164 61940 311216 61946
rect 311164 61882 311216 61888
rect 312556 60314 312584 70042
rect 318248 69556 318300 69562
rect 318248 69498 318300 69504
rect 318064 68876 318116 68882
rect 318064 68818 318116 68824
rect 316684 68808 316736 68814
rect 316684 68750 316736 68756
rect 315304 61940 315356 61946
rect 315304 61882 315356 61888
rect 313924 61396 313976 61402
rect 313924 61338 313976 61344
rect 312544 60308 312596 60314
rect 312544 60250 312596 60256
rect 313188 57248 313240 57254
rect 313188 57190 313240 57196
rect 309784 56568 309836 56574
rect 309784 56510 309836 56516
rect 307668 55888 307720 55894
rect 307668 55830 307720 55836
rect 306104 54800 306156 54806
rect 306104 54742 306156 54748
rect 309876 54800 309928 54806
rect 309876 54742 309928 54748
rect 306012 54732 306064 54738
rect 306012 54674 306064 54680
rect 309784 54732 309836 54738
rect 309784 54674 309836 54680
rect 305644 50380 305696 50386
rect 305644 50322 305696 50328
rect 305920 50380 305972 50386
rect 305920 50322 305972 50328
rect 305000 47592 305052 47598
rect 305000 47534 305052 47540
rect 305656 40730 305684 50322
rect 308496 49088 308548 49094
rect 308496 49030 308548 49036
rect 308404 46232 308456 46238
rect 308404 46174 308456 46180
rect 305644 40724 305696 40730
rect 305644 40666 305696 40672
rect 307024 40044 307076 40050
rect 307024 39986 307076 39992
rect 307036 27606 307064 39986
rect 307024 27600 307076 27606
rect 307024 27542 307076 27548
rect 306380 26376 306432 26382
rect 306380 26318 306432 26324
rect 304448 24132 304500 24138
rect 304448 24074 304500 24080
rect 304356 18760 304408 18766
rect 304356 18702 304408 18708
rect 304264 14952 304316 14958
rect 304264 14894 304316 14900
rect 304368 9110 304396 18702
rect 304460 16318 304488 24074
rect 305644 23044 305696 23050
rect 305644 22986 305696 22992
rect 305000 22840 305052 22846
rect 305000 22782 305052 22788
rect 305012 16574 305040 22782
rect 305012 16546 305592 16574
rect 304448 16312 304500 16318
rect 304448 16254 304500 16260
rect 304356 9104 304408 9110
rect 304356 9046 304408 9052
rect 305564 480 305592 16546
rect 305656 6322 305684 22986
rect 306392 22846 306420 26318
rect 307116 24880 307168 24886
rect 307116 24822 307168 24828
rect 307024 22908 307076 22914
rect 307024 22850 307076 22856
rect 306380 22840 306432 22846
rect 306380 22782 306432 22788
rect 306746 9072 306802 9081
rect 306746 9007 306802 9016
rect 305644 6316 305696 6322
rect 305644 6258 305696 6264
rect 306760 480 306788 9007
rect 307036 4010 307064 22850
rect 307128 12306 307156 24822
rect 308416 23254 308444 46174
rect 308508 43586 308536 49030
rect 309600 47592 309652 47598
rect 309600 47534 309652 47540
rect 309048 44940 309100 44946
rect 309048 44882 309100 44888
rect 308496 43580 308548 43586
rect 308496 43522 308548 43528
rect 309060 41274 309088 44882
rect 309048 41268 309100 41274
rect 309048 41210 309100 41216
rect 309612 40798 309640 47534
rect 309796 43246 309824 54674
rect 309888 43382 309916 54742
rect 312544 54664 312596 54670
rect 312544 54606 312596 54612
rect 309968 53236 310020 53242
rect 309968 53178 310020 53184
rect 309980 43518 310008 53178
rect 311164 51740 311216 51746
rect 311164 51682 311216 51688
rect 310428 50448 310480 50454
rect 310428 50390 310480 50396
rect 310440 46238 310468 50390
rect 310612 49224 310664 49230
rect 310612 49166 310664 49172
rect 310520 49156 310572 49162
rect 310520 49098 310572 49104
rect 310532 46850 310560 49098
rect 310520 46844 310572 46850
rect 310520 46786 310572 46792
rect 310624 46782 310652 49166
rect 310612 46776 310664 46782
rect 310612 46718 310664 46724
rect 310428 46232 310480 46238
rect 310428 46174 310480 46180
rect 311176 44606 311204 51682
rect 311164 44600 311216 44606
rect 311164 44542 311216 44548
rect 309968 43512 310020 43518
rect 309968 43454 310020 43460
rect 309876 43376 309928 43382
rect 309876 43318 309928 43324
rect 312268 43376 312320 43382
rect 312268 43318 312320 43324
rect 309784 43240 309836 43246
rect 309784 43182 309836 43188
rect 311900 43240 311952 43246
rect 311900 43182 311952 43188
rect 310704 41268 310756 41274
rect 310704 41210 310756 41216
rect 309600 40792 309652 40798
rect 309600 40734 309652 40740
rect 310716 36990 310744 41210
rect 311912 39846 311940 43182
rect 312280 39914 312308 43318
rect 312268 39908 312320 39914
rect 312268 39850 312320 39856
rect 311900 39840 311952 39846
rect 311900 39782 311952 39788
rect 310704 36984 310756 36990
rect 310704 36926 310756 36932
rect 311164 36644 311216 36650
rect 311164 36586 311216 36592
rect 308496 36100 308548 36106
rect 308496 36042 308548 36048
rect 308508 28966 308536 36042
rect 309784 29708 309836 29714
rect 309784 29650 309836 29656
rect 308496 28960 308548 28966
rect 308496 28902 308548 28908
rect 309796 23322 309824 29650
rect 309784 23316 309836 23322
rect 309784 23258 309836 23264
rect 308404 23248 308456 23254
rect 308404 23190 308456 23196
rect 308496 20664 308548 20670
rect 308496 20606 308548 20612
rect 307208 20392 307260 20398
rect 307208 20334 307260 20340
rect 307116 12300 307168 12306
rect 307116 12242 307168 12248
rect 307220 9654 307248 20334
rect 308404 16312 308456 16318
rect 308404 16254 308456 16260
rect 307208 9648 307260 9654
rect 307208 9590 307260 9596
rect 307942 8936 307998 8945
rect 307942 8871 307998 8880
rect 307024 4004 307076 4010
rect 307024 3946 307076 3952
rect 307956 480 307984 8871
rect 308416 2990 308444 16254
rect 308508 15094 308536 20606
rect 308496 15088 308548 15094
rect 308496 15030 308548 15036
rect 311176 11694 311204 36586
rect 312556 35222 312584 54606
rect 313200 49706 313228 57190
rect 313188 49700 313240 49706
rect 313188 49642 313240 49648
rect 313280 46844 313332 46850
rect 313280 46786 313332 46792
rect 313292 39982 313320 46786
rect 313464 46776 313516 46782
rect 313464 46718 313516 46724
rect 313476 40050 313504 46718
rect 313936 41410 313964 61338
rect 314292 56568 314344 56574
rect 314292 56510 314344 56516
rect 314304 51746 314332 56510
rect 315316 51814 315344 61882
rect 315396 60308 315448 60314
rect 315396 60250 315448 60256
rect 315408 54398 315436 60250
rect 316696 56574 316724 68750
rect 316684 56568 316736 56574
rect 316684 56510 316736 56516
rect 315396 54392 315448 54398
rect 315396 54334 315448 54340
rect 315304 51808 315356 51814
rect 315304 51750 315356 51756
rect 314292 51740 314344 51746
rect 314292 51682 314344 51688
rect 318076 48278 318104 68818
rect 318156 67176 318208 67182
rect 318156 67118 318208 67124
rect 318168 50794 318196 67118
rect 318260 61402 318288 69498
rect 320560 68678 320588 75482
rect 332600 71324 332652 71330
rect 332600 71266 332652 71272
rect 332612 68746 332640 71266
rect 334716 71256 334768 71262
rect 334716 71198 334768 71204
rect 332600 68740 332652 68746
rect 332600 68682 332652 68688
rect 320548 68672 320600 68678
rect 320548 68614 320600 68620
rect 318248 61396 318300 61402
rect 318248 61338 318300 61344
rect 334624 61396 334676 61402
rect 334624 61338 334676 61344
rect 326344 60240 326396 60246
rect 326344 60182 326396 60188
rect 322204 56568 322256 56574
rect 322204 56510 322256 56516
rect 321468 55888 321520 55894
rect 321468 55830 321520 55836
rect 319444 54528 319496 54534
rect 319444 54470 319496 54476
rect 318340 54392 318392 54398
rect 318340 54334 318392 54340
rect 318156 50788 318208 50794
rect 318156 50730 318208 50736
rect 318156 49700 318208 49706
rect 318156 49642 318208 49648
rect 318064 48272 318116 48278
rect 318064 48214 318116 48220
rect 316776 46232 316828 46238
rect 316776 46174 316828 46180
rect 313924 41404 313976 41410
rect 313924 41346 313976 41352
rect 316684 41404 316736 41410
rect 316684 41346 316736 41352
rect 313464 40044 313516 40050
rect 313464 39986 313516 39992
rect 313280 39976 313332 39982
rect 313280 39918 313332 39924
rect 315304 39432 315356 39438
rect 315304 39374 315356 39380
rect 312636 37936 312688 37942
rect 312636 37878 312688 37884
rect 312544 35216 312596 35222
rect 312544 35158 312596 35164
rect 312176 27600 312228 27606
rect 312176 27542 312228 27548
rect 312188 22370 312216 27542
rect 312648 27062 312676 37878
rect 312636 27056 312688 27062
rect 312636 26998 312688 27004
rect 315316 26042 315344 39374
rect 316592 28960 316644 28966
rect 316592 28902 316644 28908
rect 316604 28218 316632 28902
rect 316592 28212 316644 28218
rect 316592 28154 316644 28160
rect 315304 26036 315356 26042
rect 315304 25978 315356 25984
rect 312912 23316 312964 23322
rect 312912 23258 312964 23264
rect 312176 22364 312228 22370
rect 312176 22306 312228 22312
rect 312924 20330 312952 23258
rect 313280 23248 313332 23254
rect 313280 23190 313332 23196
rect 312912 20324 312964 20330
rect 312912 20266 312964 20272
rect 312544 18692 312596 18698
rect 312544 18634 312596 18640
rect 311900 12300 311952 12306
rect 311900 12242 311952 12248
rect 311164 11688 311216 11694
rect 311164 11630 311216 11636
rect 309324 9648 309376 9654
rect 309324 9590 309376 9596
rect 309336 6322 309364 9590
rect 311912 7546 311940 12242
rect 312268 9104 312320 9110
rect 312268 9046 312320 9052
rect 311900 7540 311952 7546
rect 311900 7482 311952 7488
rect 309232 6316 309284 6322
rect 309232 6258 309284 6264
rect 309324 6316 309376 6322
rect 309324 6258 309376 6264
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 308404 2984 308456 2990
rect 308404 2926 308456 2932
rect 309060 480 309088 3334
rect 309244 3194 309272 6258
rect 310244 4072 310296 4078
rect 310244 4014 310296 4020
rect 309232 3188 309284 3194
rect 309232 3130 309284 3136
rect 310256 480 310284 4014
rect 311440 2984 311492 2990
rect 311440 2926 311492 2932
rect 311452 480 311480 2926
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312280 354 312308 9046
rect 312556 7750 312584 18634
rect 312636 17672 312688 17678
rect 312636 17614 312688 17620
rect 312648 8362 312676 17614
rect 313292 16574 313320 23190
rect 315304 22364 315356 22370
rect 315304 22306 315356 22312
rect 313292 16546 313872 16574
rect 312636 8356 312688 8362
rect 312636 8298 312688 8304
rect 312544 7744 312596 7750
rect 312544 7686 312596 7692
rect 313844 480 313872 16546
rect 314752 15020 314804 15026
rect 314752 14962 314804 14968
rect 314660 11688 314712 11694
rect 314660 11630 314712 11636
rect 312606 354 312718 480
rect 312280 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 11630
rect 314764 7682 314792 14962
rect 315316 9110 315344 22306
rect 316696 11014 316724 41346
rect 316788 37942 316816 46174
rect 317328 44600 317380 44606
rect 317328 44542 317380 44548
rect 317052 43580 317104 43586
rect 317052 43522 317104 43528
rect 316776 37936 316828 37942
rect 316776 37878 316828 37884
rect 317064 37126 317092 43522
rect 317340 41342 317368 44542
rect 317328 41336 317380 41342
rect 317328 41278 317380 41284
rect 317236 40044 317288 40050
rect 317236 39986 317288 39992
rect 317052 37120 317104 37126
rect 317052 37062 317104 37068
rect 316776 36984 316828 36990
rect 316776 36926 316828 36932
rect 316788 24478 316816 36926
rect 317248 36786 317276 39986
rect 317328 39976 317380 39982
rect 317328 39918 317380 39924
rect 317340 36854 317368 39918
rect 318168 39438 318196 49642
rect 318352 48210 318380 54334
rect 318340 48204 318392 48210
rect 318340 48146 318392 48152
rect 319456 46850 319484 54470
rect 321480 53174 321508 55830
rect 321468 53168 321520 53174
rect 321468 53110 321520 53116
rect 320732 51808 320784 51814
rect 320732 51750 320784 51756
rect 319536 50380 319588 50386
rect 319536 50322 319588 50328
rect 319444 46844 319496 46850
rect 319444 46786 319496 46792
rect 319444 43512 319496 43518
rect 319444 43454 319496 43460
rect 318524 39908 318576 39914
rect 318524 39850 318576 39856
rect 318432 39840 318484 39846
rect 318432 39782 318484 39788
rect 318156 39432 318208 39438
rect 318156 39374 318208 39380
rect 318444 37262 318472 39782
rect 318432 37256 318484 37262
rect 318432 37198 318484 37204
rect 318536 37194 318564 39850
rect 318524 37188 318576 37194
rect 318524 37130 318576 37136
rect 317328 36848 317380 36854
rect 317328 36790 317380 36796
rect 316868 36780 316920 36786
rect 316868 36722 316920 36728
rect 317236 36780 317288 36786
rect 317236 36722 317288 36728
rect 316880 28966 316908 36722
rect 316868 28960 316920 28966
rect 316868 28902 316920 28908
rect 318064 28212 318116 28218
rect 318064 28154 318116 28160
rect 316776 24472 316828 24478
rect 316776 24414 316828 24420
rect 316684 11008 316736 11014
rect 316684 10950 316736 10956
rect 318076 10946 318104 28154
rect 319456 13870 319484 43454
rect 319548 42090 319576 50322
rect 320744 46238 320772 51750
rect 320824 51740 320876 51746
rect 320824 51682 320876 51688
rect 320732 46232 320784 46238
rect 320732 46174 320784 46180
rect 320836 44334 320864 51682
rect 321008 48204 321060 48210
rect 321008 48146 321060 48152
rect 320824 44328 320876 44334
rect 320824 44270 320876 44276
rect 319536 42084 319588 42090
rect 319536 42026 319588 42032
rect 320824 37256 320876 37262
rect 320824 37198 320876 37204
rect 319628 28960 319680 28966
rect 319628 28902 319680 28908
rect 319536 24472 319588 24478
rect 319536 24414 319588 24420
rect 319444 13864 319496 13870
rect 319444 13806 319496 13812
rect 319444 11008 319496 11014
rect 319444 10950 319496 10956
rect 318064 10940 318116 10946
rect 318064 10882 318116 10888
rect 315304 9104 315356 9110
rect 315304 9046 315356 9052
rect 316224 8356 316276 8362
rect 316224 8298 316276 8304
rect 314752 7676 314804 7682
rect 314752 7618 314804 7624
rect 316236 480 316264 8298
rect 317420 7540 317472 7546
rect 317420 7482 317472 7488
rect 317432 3942 317460 7482
rect 318524 4004 318576 4010
rect 318524 3946 318576 3952
rect 317420 3936 317472 3942
rect 317420 3878 317472 3884
rect 317328 3188 317380 3194
rect 317328 3130 317380 3136
rect 317340 480 317368 3130
rect 318536 480 318564 3946
rect 319456 3482 319484 10950
rect 319548 5574 319576 24414
rect 319640 12102 319668 28902
rect 320088 27056 320140 27062
rect 320088 26998 320140 27004
rect 320100 24206 320128 26998
rect 320180 26036 320232 26042
rect 320180 25978 320232 25984
rect 320088 24200 320140 24206
rect 320088 24142 320140 24148
rect 320192 16574 320220 25978
rect 320192 16546 320496 16574
rect 319812 15088 319864 15094
rect 319812 15030 319864 15036
rect 319628 12096 319680 12102
rect 319628 12038 319680 12044
rect 319536 5568 319588 5574
rect 319536 5510 319588 5516
rect 319456 3454 319760 3482
rect 319732 480 319760 3454
rect 319824 3330 319852 15030
rect 319812 3324 319864 3330
rect 319812 3266 319864 3272
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 320732 14952 320784 14958
rect 320732 14894 320784 14900
rect 320744 12170 320772 14894
rect 320732 12164 320784 12170
rect 320732 12106 320784 12112
rect 320836 9586 320864 37198
rect 320916 37188 320968 37194
rect 320916 37130 320968 37136
rect 320928 9654 320956 37130
rect 321020 24886 321048 48146
rect 322216 41614 322244 56510
rect 323768 54596 323820 54602
rect 323768 54538 323820 54544
rect 323676 50788 323728 50794
rect 323676 50730 323728 50736
rect 323584 48272 323636 48278
rect 323584 48214 323636 48220
rect 322848 46844 322900 46850
rect 322848 46786 322900 46792
rect 322204 41608 322256 41614
rect 322204 41550 322256 41556
rect 322860 41410 322888 46786
rect 323032 44328 323084 44334
rect 323032 44270 323084 44276
rect 322848 41404 322900 41410
rect 322848 41346 322900 41352
rect 321100 40792 321152 40798
rect 321100 40734 321152 40740
rect 321112 26042 321140 40734
rect 322940 40724 322992 40730
rect 322940 40666 322992 40672
rect 322952 37670 322980 40666
rect 322940 37664 322992 37670
rect 322940 37606 322992 37612
rect 322756 37120 322808 37126
rect 322756 37062 322808 37068
rect 322768 29714 322796 37062
rect 323044 36650 323072 44270
rect 323032 36644 323084 36650
rect 323032 36586 323084 36592
rect 323596 31754 323624 48214
rect 323688 34474 323716 50730
rect 323780 43518 323808 54538
rect 326356 53106 326384 60182
rect 330484 53168 330536 53174
rect 330484 53110 330536 53116
rect 326344 53100 326396 53106
rect 326344 53042 326396 53048
rect 330496 50862 330524 53110
rect 330484 50856 330536 50862
rect 330484 50798 330536 50804
rect 323768 43512 323820 43518
rect 323768 43454 323820 43460
rect 326068 43512 326120 43518
rect 326068 43454 326120 43460
rect 324964 41608 325016 41614
rect 324964 41550 325016 41556
rect 323768 36712 323820 36718
rect 323768 36654 323820 36660
rect 323676 34468 323728 34474
rect 323676 34410 323728 34416
rect 323584 31748 323636 31754
rect 323584 31690 323636 31696
rect 322756 29708 322808 29714
rect 322756 29650 322808 29656
rect 323780 27062 323808 36654
rect 324320 35216 324372 35222
rect 324320 35158 324372 35164
rect 323768 27056 323820 27062
rect 323768 26998 323820 27004
rect 324332 26994 324360 35158
rect 324976 27674 325004 41550
rect 325056 41336 325108 41342
rect 325056 41278 325108 41284
rect 325068 30326 325096 41278
rect 326080 36718 326108 43454
rect 334636 42158 334664 61338
rect 334728 59362 334756 71198
rect 336752 69018 336780 76638
rect 361580 76628 361632 76634
rect 361580 76570 361632 76576
rect 347780 72616 347832 72622
rect 347780 72558 347832 72564
rect 345664 71188 345716 71194
rect 345664 71130 345716 71136
rect 336740 69012 336792 69018
rect 336740 68954 336792 68960
rect 339500 69012 339552 69018
rect 339500 68954 339552 68960
rect 339512 65822 339540 68954
rect 340144 68740 340196 68746
rect 340144 68682 340196 68688
rect 339500 65816 339552 65822
rect 339500 65758 339552 65764
rect 340156 61742 340184 68682
rect 340144 61736 340196 61742
rect 340144 61678 340196 61684
rect 344284 61736 344336 61742
rect 344284 61678 344336 61684
rect 334716 59356 334768 59362
rect 334716 59298 334768 59304
rect 337384 59356 337436 59362
rect 337384 59298 337436 59304
rect 336096 50856 336148 50862
rect 336096 50798 336148 50804
rect 334624 42152 334676 42158
rect 334624 42094 334676 42100
rect 327724 41404 327776 41410
rect 327724 41346 327776 41352
rect 327080 37936 327132 37942
rect 327080 37878 327132 37884
rect 326160 37664 326212 37670
rect 326160 37606 326212 37612
rect 326068 36712 326120 36718
rect 326068 36654 326120 36660
rect 326172 34950 326200 37606
rect 326160 34944 326212 34950
rect 326160 34886 326212 34892
rect 326344 31748 326396 31754
rect 326344 31690 326396 31696
rect 325056 30320 325108 30326
rect 325056 30262 325108 30268
rect 324964 27668 325016 27674
rect 324964 27610 325016 27616
rect 321192 26988 321244 26994
rect 321192 26930 321244 26936
rect 324320 26988 324372 26994
rect 324320 26930 324372 26936
rect 321100 26036 321152 26042
rect 321100 25978 321152 25984
rect 321008 24880 321060 24886
rect 321008 24822 321060 24828
rect 321204 13802 321232 26930
rect 323584 24880 323636 24886
rect 323584 24822 323636 24828
rect 323596 15978 323624 24822
rect 324964 24200 325016 24206
rect 324964 24142 325016 24148
rect 323584 15972 323636 15978
rect 323584 15914 323636 15920
rect 324976 14958 325004 24142
rect 326356 24138 326384 31690
rect 327092 31006 327120 37878
rect 327080 31000 327132 31006
rect 327080 30942 327132 30948
rect 327080 27668 327132 27674
rect 327080 27610 327132 27616
rect 326344 24132 326396 24138
rect 326344 24074 326396 24080
rect 327092 21690 327120 27610
rect 327080 21684 327132 21690
rect 327080 21626 327132 21632
rect 327080 20324 327132 20330
rect 327080 20266 327132 20272
rect 327092 16574 327120 20266
rect 327092 16546 327212 16574
rect 324964 14952 325016 14958
rect 324964 14894 325016 14900
rect 322204 13864 322256 13870
rect 322204 13806 322256 13812
rect 321192 13796 321244 13802
rect 321192 13738 321244 13744
rect 320916 9648 320968 9654
rect 320916 9590 320968 9596
rect 320824 9580 320876 9586
rect 320824 9522 320876 9528
rect 322112 3324 322164 3330
rect 322112 3266 322164 3272
rect 322124 480 322152 3266
rect 322216 3262 322244 13806
rect 326344 13796 326396 13802
rect 326344 13738 326396 13744
rect 322296 12096 322348 12102
rect 322296 12038 322348 12044
rect 322308 3398 322336 12038
rect 322388 10940 322440 10946
rect 322388 10882 322440 10888
rect 322400 4010 322428 10882
rect 324688 9648 324740 9654
rect 324688 9590 324740 9596
rect 323308 7744 323360 7750
rect 323308 7686 323360 7692
rect 322388 4004 322440 4010
rect 322388 3946 322440 3952
rect 322296 3392 322348 3398
rect 322296 3334 322348 3340
rect 322204 3256 322256 3262
rect 322204 3198 322256 3204
rect 323320 480 323348 7686
rect 324700 6526 324728 9590
rect 324780 9580 324832 9586
rect 324780 9522 324832 9528
rect 324688 6520 324740 6526
rect 324688 6462 324740 6468
rect 324792 6458 324820 9522
rect 324780 6452 324832 6458
rect 324780 6394 324832 6400
rect 326356 5574 326384 13738
rect 327080 7676 327132 7682
rect 327080 7618 327132 7624
rect 324412 5568 324464 5574
rect 324412 5510 324464 5516
rect 326344 5568 326396 5574
rect 326344 5510 326396 5516
rect 324424 480 324452 5510
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 325620 480 325648 3334
rect 326804 3256 326856 3262
rect 326804 3198 326856 3204
rect 326816 480 326844 3198
rect 327092 3126 327120 7618
rect 327184 6914 327212 16546
rect 327736 11694 327764 41346
rect 330484 36848 330536 36854
rect 330484 36790 330536 36796
rect 329196 34468 329248 34474
rect 329196 34410 329248 34416
rect 327908 30320 327960 30326
rect 327908 30262 327960 30268
rect 327920 24206 327948 30262
rect 329104 27056 329156 27062
rect 329104 26998 329156 27004
rect 329012 26036 329064 26042
rect 329012 25978 329064 25984
rect 327908 24200 327960 24206
rect 327908 24142 327960 24148
rect 329024 22710 329052 25978
rect 329012 22704 329064 22710
rect 329012 22646 329064 22652
rect 329116 13258 329144 26998
rect 329208 21758 329236 34410
rect 329196 21752 329248 21758
rect 329196 21694 329248 21700
rect 330496 18698 330524 36790
rect 330576 36780 330628 36786
rect 330576 36722 330628 36728
rect 330588 18834 330616 36722
rect 336004 36712 336056 36718
rect 336004 36654 336056 36660
rect 333244 34944 333296 34950
rect 333244 34886 333296 34892
rect 330668 31000 330720 31006
rect 330668 30942 330720 30948
rect 330680 19310 330708 30942
rect 333256 26042 333284 34886
rect 334624 26988 334676 26994
rect 334624 26930 334676 26936
rect 333244 26036 333296 26042
rect 333244 25978 333296 25984
rect 330668 19304 330720 19310
rect 330668 19246 330720 19252
rect 330576 18828 330628 18834
rect 330576 18770 330628 18776
rect 330484 18692 330536 18698
rect 330484 18634 330536 18640
rect 333244 15972 333296 15978
rect 333244 15914 333296 15920
rect 329104 13252 329156 13258
rect 329104 13194 329156 13200
rect 329104 12096 329156 12102
rect 329104 12038 329156 12044
rect 327724 11688 327776 11694
rect 327724 11630 327776 11636
rect 327184 6886 328040 6914
rect 327080 3120 327132 3126
rect 327080 3062 327132 3068
rect 328012 480 328040 6886
rect 329116 3398 329144 12038
rect 330484 11688 330536 11694
rect 330484 11630 330536 11636
rect 329196 4004 329248 4010
rect 329196 3946 329248 3952
rect 329104 3392 329156 3398
rect 329104 3334 329156 3340
rect 329208 480 329236 3946
rect 330392 3936 330444 3942
rect 330392 3878 330444 3884
rect 330404 480 330432 3878
rect 330496 3058 330524 11630
rect 330760 9104 330812 9110
rect 330760 9046 330812 9052
rect 330772 6390 330800 9046
rect 333256 6594 333284 15914
rect 334636 15026 334664 26930
rect 334808 22704 334860 22710
rect 334808 22646 334860 22652
rect 334716 19304 334768 19310
rect 334716 19246 334768 19252
rect 334624 15020 334676 15026
rect 334624 14962 334676 14968
rect 334624 13252 334676 13258
rect 334624 13194 334676 13200
rect 333244 6588 333296 6594
rect 333244 6530 333296 6536
rect 334072 6520 334124 6526
rect 334072 6462 334124 6468
rect 333980 6452 334032 6458
rect 333980 6394 334032 6400
rect 330760 6384 330812 6390
rect 330760 6326 330812 6332
rect 332692 5568 332744 5574
rect 332692 5510 332744 5516
rect 331588 3120 331640 3126
rect 331588 3062 331640 3068
rect 330484 3052 330536 3058
rect 330484 2994 330536 3000
rect 331600 480 331628 3062
rect 332704 480 332732 5510
rect 333992 3942 334020 6394
rect 333980 3936 334032 3942
rect 333980 3878 334032 3884
rect 334084 3330 334112 6462
rect 334072 3324 334124 3330
rect 334072 3266 334124 3272
rect 333888 3052 333940 3058
rect 333888 2994 333940 3000
rect 333900 480 333928 2994
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 13194
rect 334728 7682 334756 19246
rect 334820 15978 334848 22646
rect 334808 15972 334860 15978
rect 334808 15914 334860 15920
rect 336016 9654 336044 36654
rect 336108 28966 336136 50798
rect 336188 42084 336240 42090
rect 336188 42026 336240 42032
rect 336200 31890 336228 42026
rect 337396 33182 337424 59298
rect 338764 46232 338816 46238
rect 338764 46174 338816 46180
rect 337936 39432 337988 39438
rect 337936 39374 337988 39380
rect 337948 37262 337976 39374
rect 338776 38486 338804 46174
rect 340144 42152 340196 42158
rect 340144 42094 340196 42100
rect 338764 38480 338816 38486
rect 338764 38422 338816 38428
rect 337936 37256 337988 37262
rect 337936 37198 337988 37204
rect 337384 33176 337436 33182
rect 337384 33118 337436 33124
rect 339960 33176 340012 33182
rect 339960 33118 340012 33124
rect 336188 31884 336240 31890
rect 336188 31826 336240 31832
rect 339972 30326 340000 33118
rect 340156 33114 340184 42094
rect 340788 37256 340840 37262
rect 340788 37198 340840 37204
rect 340696 36644 340748 36650
rect 340696 36586 340748 36592
rect 340144 33108 340196 33114
rect 340144 33050 340196 33056
rect 340708 33046 340736 36586
rect 340800 34474 340828 37198
rect 340788 34468 340840 34474
rect 340788 34410 340840 34416
rect 340696 33040 340748 33046
rect 340696 32982 340748 32988
rect 343640 33040 343692 33046
rect 343640 32982 343692 32988
rect 342904 31884 342956 31890
rect 342904 31826 342956 31832
rect 339960 30320 340012 30326
rect 339960 30262 340012 30268
rect 336096 28960 336148 28966
rect 336096 28902 336148 28908
rect 341064 28960 341116 28966
rect 341064 28902 341116 28908
rect 341076 22846 341104 28902
rect 342260 24132 342312 24138
rect 342260 24074 342312 24080
rect 340052 22840 340104 22846
rect 340052 22782 340104 22788
rect 341064 22840 341116 22846
rect 341064 22782 341116 22788
rect 338764 18828 338816 18834
rect 338764 18770 338816 18776
rect 336004 9648 336056 9654
rect 336004 9590 336056 9596
rect 338776 9110 338804 18770
rect 339316 18692 339368 18698
rect 339316 18634 339368 18640
rect 339040 15972 339092 15978
rect 339040 15914 339092 15920
rect 339052 11014 339080 15914
rect 339328 15094 339356 18634
rect 339316 15088 339368 15094
rect 339316 15030 339368 15036
rect 340064 12510 340092 22782
rect 341524 21752 341576 21758
rect 341524 21694 341576 21700
rect 340144 21684 340196 21690
rect 340144 21626 340196 21632
rect 340156 18698 340184 21626
rect 340144 18692 340196 18698
rect 340144 18634 340196 18640
rect 340236 15020 340288 15026
rect 340236 14962 340288 14968
rect 340052 12504 340104 12510
rect 340052 12446 340104 12452
rect 339040 11008 339092 11014
rect 339040 10950 339092 10956
rect 338764 9104 338816 9110
rect 338764 9046 338816 9052
rect 334716 7676 334768 7682
rect 334716 7618 334768 7624
rect 338672 6588 338724 6594
rect 338672 6530 338724 6536
rect 336280 3392 336332 3398
rect 336280 3334 336332 3340
rect 336292 480 336320 3334
rect 337476 3324 337528 3330
rect 337476 3266 337528 3272
rect 337488 480 337516 3266
rect 338684 480 338712 6530
rect 340248 6458 340276 14962
rect 341536 13734 341564 21694
rect 342272 16862 342300 24074
rect 342260 16856 342312 16862
rect 342260 16798 342312 16804
rect 342916 15978 342944 31826
rect 343652 30258 343680 32982
rect 343640 30252 343692 30258
rect 343640 30194 343692 30200
rect 343640 26036 343692 26042
rect 343640 25978 343692 25984
rect 343652 16574 343680 25978
rect 344296 21690 344324 61678
rect 345676 37262 345704 71130
rect 345756 65816 345808 65822
rect 345756 65758 345808 65764
rect 345768 51406 345796 65758
rect 345756 51400 345808 51406
rect 345756 51342 345808 51348
rect 347136 38480 347188 38486
rect 347136 38422 347188 38428
rect 345664 37256 345716 37262
rect 345664 37198 345716 37204
rect 345940 33108 345992 33114
rect 345940 33050 345992 33056
rect 345020 30320 345072 30326
rect 345020 30262 345072 30268
rect 344468 29708 344520 29714
rect 344468 29650 344520 29656
rect 344376 24200 344428 24206
rect 344376 24142 344428 24148
rect 344284 21684 344336 21690
rect 344284 21626 344336 21632
rect 343652 16546 344324 16574
rect 342904 15972 342956 15978
rect 342904 15914 342956 15920
rect 342812 15088 342864 15094
rect 342812 15030 342864 15036
rect 341524 13728 341576 13734
rect 341524 13670 341576 13676
rect 342720 11008 342772 11014
rect 342720 10950 342772 10956
rect 342168 9648 342220 9654
rect 342168 9590 342220 9596
rect 340236 6452 340288 6458
rect 340236 6394 340288 6400
rect 339868 6316 339920 6322
rect 339868 6258 339920 6264
rect 339880 480 339908 6258
rect 340972 3936 341024 3942
rect 340972 3878 341024 3884
rect 340984 480 341012 3878
rect 342180 480 342208 9590
rect 342732 490 342760 10950
rect 342824 3942 342852 15030
rect 342996 12504 343048 12510
rect 342996 12446 343048 12452
rect 343008 6322 343036 12446
rect 343640 6384 343692 6390
rect 343640 6326 343692 6332
rect 342996 6316 343048 6322
rect 342996 6258 343048 6264
rect 343652 4146 343680 6326
rect 343640 4140 343692 4146
rect 343640 4082 343692 4088
rect 342812 3936 342864 3942
rect 342812 3878 342864 3884
rect 344296 3482 344324 16546
rect 344388 4078 344416 24142
rect 344480 24138 344508 29650
rect 344468 24132 344520 24138
rect 344468 24074 344520 24080
rect 345032 16574 345060 30262
rect 345952 28218 345980 33050
rect 347044 30252 347096 30258
rect 347044 30194 347096 30200
rect 345940 28212 345992 28218
rect 345940 28154 345992 28160
rect 347056 20670 347084 30194
rect 347148 28966 347176 38422
rect 347136 28960 347188 28966
rect 347136 28902 347188 28908
rect 347044 20664 347096 20670
rect 347044 20606 347096 20612
rect 346400 16856 346452 16862
rect 346400 16798 346452 16804
rect 346412 16574 346440 16798
rect 347792 16574 347820 72558
rect 349068 72548 349120 72554
rect 349068 72490 349120 72496
rect 348700 66972 348752 66978
rect 348700 66914 348752 66920
rect 348712 62830 348740 66914
rect 349080 65618 349108 72490
rect 349804 69896 349856 69902
rect 349804 69838 349856 69844
rect 349068 65612 349120 65618
rect 349068 65554 349120 65560
rect 348700 62824 348752 62830
rect 348700 62766 348752 62772
rect 348424 51400 348476 51406
rect 348424 51342 348476 51348
rect 345032 16546 345336 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 344376 4072 344428 4078
rect 344376 4014 344428 4020
rect 344296 3454 344600 3482
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342732 462 342944 490
rect 344572 480 344600 3454
rect 342916 354 342944 462
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346964 480 346992 16546
rect 347872 15972 347924 15978
rect 347872 15914 347924 15920
rect 347136 14952 347188 14958
rect 347136 14894 347188 14900
rect 347044 13728 347096 13734
rect 347044 13670 347096 13676
rect 347056 3126 347084 13670
rect 347148 11014 347176 14894
rect 347884 12102 347912 15914
rect 347872 12096 347924 12102
rect 347872 12038 347924 12044
rect 347136 11008 347188 11014
rect 347136 10950 347188 10956
rect 347044 3120 347096 3126
rect 347044 3062 347096 3068
rect 348068 480 348096 16546
rect 348436 14414 348464 51342
rect 348516 37256 348568 37262
rect 348516 37198 348568 37204
rect 348528 27606 348556 37198
rect 348516 27600 348568 27606
rect 348516 27542 348568 27548
rect 349816 26042 349844 69838
rect 359556 68672 359608 68678
rect 359556 68614 359608 68620
rect 359464 65612 359516 65618
rect 359464 65554 359516 65560
rect 351920 62824 351972 62830
rect 351920 62766 351972 62772
rect 351932 58818 351960 62766
rect 351920 58812 351972 58818
rect 351920 58754 351972 58760
rect 350540 53100 350592 53106
rect 350540 53042 350592 53048
rect 350552 46238 350580 53042
rect 350540 46232 350592 46238
rect 350540 46174 350592 46180
rect 359476 43790 359504 65554
rect 359568 61470 359596 68614
rect 359556 61464 359608 61470
rect 359556 61406 359608 61412
rect 359464 43784 359516 43790
rect 359464 43726 359516 43732
rect 353944 34468 353996 34474
rect 353944 34410 353996 34416
rect 352564 28960 352616 28966
rect 352564 28902 352616 28908
rect 349804 26036 349856 26042
rect 349804 25978 349856 25984
rect 349896 24132 349948 24138
rect 349896 24074 349948 24080
rect 349908 20670 349936 24074
rect 349804 20664 349856 20670
rect 349804 20606 349856 20612
rect 349896 20664 349948 20670
rect 349896 20606 349948 20612
rect 349160 18692 349212 18698
rect 349160 18634 349212 18640
rect 348424 14408 348476 14414
rect 348424 14350 348476 14356
rect 349172 3398 349200 18634
rect 349816 15774 349844 20606
rect 349804 15768 349856 15774
rect 349804 15710 349856 15716
rect 352288 15768 352340 15774
rect 352288 15710 352340 15716
rect 350908 14408 350960 14414
rect 350908 14350 350960 14356
rect 349252 11008 349304 11014
rect 349252 10950 349304 10956
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 349264 480 349292 10950
rect 350920 10402 350948 14350
rect 350908 10396 350960 10402
rect 350908 10338 350960 10344
rect 352300 9178 352328 15710
rect 352288 9172 352340 9178
rect 352288 9114 352340 9120
rect 351460 9104 351512 9110
rect 351460 9046 351512 9052
rect 351472 5914 351500 9046
rect 351460 5908 351512 5914
rect 351460 5850 351512 5856
rect 352576 4146 352604 28902
rect 353300 28212 353352 28218
rect 353300 28154 353352 28160
rect 352656 27600 352708 27606
rect 352656 27542 352708 27548
rect 352668 22098 352696 27542
rect 353312 24138 353340 28154
rect 353300 24132 353352 24138
rect 353300 24074 353352 24080
rect 352656 22092 352708 22098
rect 352656 22034 352708 22040
rect 352656 21684 352708 21690
rect 352656 21626 352708 21632
rect 352668 12170 352696 21626
rect 353956 13802 353984 34410
rect 360200 34400 360252 34406
rect 360200 34342 360252 34348
rect 359280 24132 359332 24138
rect 359280 24074 359332 24080
rect 358084 22840 358136 22846
rect 358084 22782 358136 22788
rect 357164 22092 357216 22098
rect 357164 22034 357216 22040
rect 355600 20664 355652 20670
rect 355600 20606 355652 20612
rect 355612 17678 355640 20606
rect 357176 18698 357204 22034
rect 357164 18692 357216 18698
rect 357164 18634 357216 18640
rect 355600 17672 355652 17678
rect 355600 17614 355652 17620
rect 353944 13796 353996 13802
rect 353944 13738 353996 13744
rect 356704 13796 356756 13802
rect 356704 13738 356756 13744
rect 352656 12164 352708 12170
rect 352656 12106 352708 12112
rect 356336 7676 356388 7682
rect 356336 7618 356388 7624
rect 352840 6452 352892 6458
rect 352840 6394 352892 6400
rect 351644 4140 351696 4146
rect 351644 4082 351696 4088
rect 352564 4140 352616 4146
rect 352564 4082 352616 4088
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 351656 480 351684 4082
rect 352852 480 352880 6394
rect 353300 5908 353352 5914
rect 353300 5850 353352 5856
rect 353312 4010 353340 5850
rect 355232 4140 355284 4146
rect 355232 4082 355284 4088
rect 353300 4004 353352 4010
rect 353300 3946 353352 3952
rect 354036 3120 354088 3126
rect 354036 3062 354088 3068
rect 354048 480 354076 3062
rect 355244 480 355272 4082
rect 356348 480 356376 7618
rect 356716 5982 356744 13738
rect 358096 12442 358124 22782
rect 359292 20670 359320 24074
rect 359280 20664 359332 20670
rect 359280 20606 359332 20612
rect 360212 16574 360240 34342
rect 361592 16574 361620 76570
rect 398840 76560 398892 76566
rect 398840 76502 398892 76508
rect 396078 71360 396134 71369
rect 396078 71295 396134 71304
rect 380900 64252 380952 64258
rect 380900 64194 380952 64200
rect 361672 61464 361724 61470
rect 361672 61406 361724 61412
rect 361684 55894 361712 61406
rect 369124 58812 369176 58818
rect 369124 58754 369176 58760
rect 361672 55888 361724 55894
rect 361672 55830 361724 55836
rect 362224 46232 362276 46238
rect 362224 46174 362276 46180
rect 362236 36650 362264 46174
rect 363604 43784 363656 43790
rect 363604 43726 363656 43732
rect 362224 36644 362276 36650
rect 362224 36586 362276 36592
rect 363616 26110 363644 43726
rect 367744 36644 367796 36650
rect 367744 36586 367796 36592
rect 363604 26104 363656 26110
rect 363604 26046 363656 26052
rect 367560 26104 367612 26110
rect 367560 26046 367612 26052
rect 364984 26036 365036 26042
rect 364984 25978 365036 25984
rect 360212 16546 361160 16574
rect 361592 16546 361896 16574
rect 358084 12436 358136 12442
rect 358084 12378 358136 12384
rect 357532 12164 357584 12170
rect 357532 12106 357584 12112
rect 357164 6316 357216 6322
rect 357164 6258 357216 6264
rect 356704 5976 356756 5982
rect 356704 5918 356756 5924
rect 357176 4146 357204 6258
rect 357164 4140 357216 4146
rect 357164 4082 357216 4088
rect 357544 480 357572 12106
rect 359464 12096 359516 12102
rect 359464 12038 359516 12044
rect 358728 4072 358780 4078
rect 358728 4014 358780 4020
rect 358740 480 358768 4014
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 12038
rect 361132 480 361160 16546
rect 361580 12436 361632 12442
rect 361580 12378 361632 12384
rect 361592 9110 361620 12378
rect 361580 9104 361632 9110
rect 361580 9046 361632 9052
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 364996 13938 365024 25978
rect 367572 20670 367600 26046
rect 365076 20664 365128 20670
rect 365076 20606 365128 20612
rect 367560 20664 367612 20670
rect 367560 20606 367612 20612
rect 365088 15026 365116 20606
rect 367756 17678 367784 36586
rect 369136 32570 369164 58754
rect 377404 55888 377456 55894
rect 377404 55830 377456 55836
rect 377416 35358 377444 55830
rect 377404 35352 377456 35358
rect 377404 35294 377456 35300
rect 369124 32564 369176 32570
rect 369124 32506 369176 32512
rect 379520 32564 379572 32570
rect 379520 32506 379572 32512
rect 379532 28966 379560 32506
rect 379520 28960 379572 28966
rect 379520 28902 379572 28908
rect 375380 28892 375432 28898
rect 375380 28834 375432 28840
rect 368480 25968 368532 25974
rect 368480 25910 368532 25916
rect 365720 17672 365772 17678
rect 365720 17614 365772 17620
rect 367744 17672 367796 17678
rect 367744 17614 367796 17620
rect 365076 15020 365128 15026
rect 365076 14962 365128 14968
rect 364984 13932 365036 13938
rect 364984 13874 365036 13880
rect 365732 10402 365760 17614
rect 368492 16574 368520 25910
rect 371240 20664 371292 20670
rect 371240 20606 371292 20612
rect 369124 18692 369176 18698
rect 369124 18634 369176 18640
rect 368492 16546 369072 16574
rect 367744 13932 367796 13938
rect 367744 13874 367796 13880
rect 363512 10396 363564 10402
rect 363512 10338 363564 10344
rect 365720 10396 365772 10402
rect 365720 10338 365772 10344
rect 362960 5976 363012 5982
rect 362960 5918 363012 5924
rect 362972 3058 363000 5918
rect 362960 3052 363012 3058
rect 362960 2994 363012 3000
rect 363524 480 363552 10338
rect 364616 9172 364668 9178
rect 364616 9114 364668 9120
rect 364628 480 364656 9114
rect 367008 4140 367060 4146
rect 367008 4082 367060 4088
rect 365812 3052 365864 3058
rect 365812 2994 365864 3000
rect 365824 480 365852 2994
rect 367020 480 367048 4082
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 13874
rect 369044 3482 369072 16546
rect 369136 3942 369164 18634
rect 370504 15020 370556 15026
rect 370504 14962 370556 14968
rect 370516 4010 370544 14962
rect 370228 4004 370280 4010
rect 370228 3946 370280 3952
rect 370504 4004 370556 4010
rect 370504 3946 370556 3952
rect 369124 3936 369176 3942
rect 369124 3878 369176 3884
rect 369044 3454 369440 3482
rect 369412 480 369440 3454
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370240 354 370268 3946
rect 370566 354 370678 480
rect 370240 326 370678 354
rect 371252 354 371280 20606
rect 375392 16574 375420 28834
rect 377404 17672 377456 17678
rect 377404 17614 377456 17620
rect 375392 16546 376064 16574
rect 374092 10396 374144 10402
rect 374092 10338 374144 10344
rect 374000 4072 374052 4078
rect 374000 4014 374052 4020
rect 372896 3936 372948 3942
rect 372896 3878 372948 3884
rect 372908 480 372936 3878
rect 374012 2122 374040 4014
rect 374104 3398 374132 10338
rect 374092 3392 374144 3398
rect 374092 3334 374144 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374012 2094 374132 2122
rect 374104 480 374132 2094
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377416 8294 377444 17614
rect 380912 16574 380940 64194
rect 394698 48920 394754 48929
rect 394698 48855 394754 48864
rect 381544 35352 381596 35358
rect 381544 35294 381596 35300
rect 381556 23458 381584 35294
rect 382280 31612 382332 31618
rect 382280 31554 382332 31560
rect 381544 23452 381596 23458
rect 381544 23394 381596 23400
rect 380912 16546 381216 16574
rect 377680 9104 377732 9110
rect 377680 9046 377732 9052
rect 377404 8288 377456 8294
rect 377404 8230 377456 8236
rect 377692 480 377720 9046
rect 379980 8288 380032 8294
rect 379980 8230 380032 8236
rect 378876 4004 378928 4010
rect 378876 3946 378928 3952
rect 378888 480 378916 3946
rect 379992 480 380020 8230
rect 381188 480 381216 16546
rect 382292 3210 382320 31554
rect 389180 31544 389232 31550
rect 389180 31486 389232 31492
rect 382924 28960 382976 28966
rect 382924 28902 382976 28908
rect 382936 12034 382964 28902
rect 385040 26920 385092 26926
rect 385040 26862 385092 26868
rect 384304 23452 384356 23458
rect 384304 23394 384356 23400
rect 384316 16574 384344 23394
rect 385052 16574 385080 26862
rect 389192 16574 389220 31486
rect 390560 25900 390612 25906
rect 390560 25842 390612 25848
rect 384316 16546 384436 16574
rect 385052 16546 386000 16574
rect 389192 16546 389496 16574
rect 384304 14884 384356 14890
rect 384304 14826 384356 14832
rect 382372 12028 382424 12034
rect 382372 11970 382424 11976
rect 382924 12028 382976 12034
rect 382924 11970 382976 11976
rect 382384 3398 382412 11970
rect 382372 3392 382424 3398
rect 382372 3334 382424 3340
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 382292 3182 382412 3210
rect 382384 480 382412 3182
rect 383580 480 383608 3334
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 14826
rect 384408 3262 384436 16546
rect 384396 3256 384448 3262
rect 384396 3198 384448 3204
rect 385972 480 386000 16546
rect 387800 14816 387852 14822
rect 387800 14758 387852 14764
rect 387156 3256 387208 3262
rect 387156 3198 387208 3204
rect 387168 480 387196 3198
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 387812 354 387840 14758
rect 389468 480 389496 16546
rect 389824 12028 389876 12034
rect 389824 11970 389876 11976
rect 389836 4146 389864 11970
rect 389824 4140 389876 4146
rect 389824 4082 389876 4088
rect 390572 3210 390600 25842
rect 394712 16574 394740 48855
rect 394712 16546 395384 16574
rect 390652 14748 390704 14754
rect 390652 14690 390704 14696
rect 390664 3398 390692 14690
rect 392582 10296 392638 10305
rect 392582 10231 392638 10240
rect 390652 3392 390704 3398
rect 390652 3334 390704 3340
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 390572 3182 390692 3210
rect 390664 480 390692 3182
rect 391860 480 391888 3334
rect 388230 354 388342 480
rect 387812 326 388342 354
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 10231
rect 394240 4140 394292 4146
rect 394240 4082 394292 4088
rect 394252 480 394280 4082
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 71295
rect 397460 28824 397512 28830
rect 397460 28766 397512 28772
rect 397472 16574 397500 28766
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3210 398880 76502
rect 407120 68604 407172 68610
rect 407120 68546 407172 68552
rect 407132 66230 407160 68546
rect 407120 66224 407172 66230
rect 407120 66166 407172 66172
rect 410524 66224 410576 66230
rect 410524 66166 410576 66172
rect 410536 54126 410564 66166
rect 410524 54120 410576 54126
rect 410524 54062 410576 54068
rect 413928 54120 413980 54126
rect 413928 54062 413980 54068
rect 413940 49706 413968 54062
rect 413928 49700 413980 49706
rect 413928 49642 413980 49648
rect 404360 36576 404412 36582
rect 404360 36518 404412 36524
rect 402980 20256 403032 20262
rect 402980 20198 403032 20204
rect 398932 17604 398984 17610
rect 398932 17546 398984 17552
rect 398944 3398 398972 17546
rect 402992 16574 403020 20198
rect 402992 16546 403664 16574
rect 400864 14680 400916 14686
rect 400864 14622 400916 14628
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 14622
rect 402520 11960 402572 11966
rect 402520 11902 402572 11908
rect 402532 480 402560 11902
rect 403636 480 403664 16546
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 36518
rect 407120 28756 407172 28762
rect 407120 28698 407172 28704
rect 406016 11892 406068 11898
rect 406016 11834 406068 11840
rect 406028 480 406056 11834
rect 407132 1834 407160 28698
rect 409878 20224 409934 20233
rect 409878 20159 409934 20168
rect 409892 16574 409920 20159
rect 414018 20088 414074 20097
rect 414018 20023 414074 20032
rect 414032 16574 414060 20023
rect 409892 16546 410840 16574
rect 414032 16546 414336 16574
rect 409142 11792 409198 11801
rect 409142 11727 409198 11736
rect 407212 9036 407264 9042
rect 407212 8978 407264 8984
rect 407120 1828 407172 1834
rect 407120 1770 407172 1776
rect 407224 480 407252 8978
rect 408408 1828 408460 1834
rect 408408 1770 408460 1776
rect 408420 480 408448 1770
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 11727
rect 410812 480 410840 16546
rect 411904 15904 411956 15910
rect 411904 15846 411956 15852
rect 411916 480 411944 15846
rect 412638 11656 412694 11665
rect 412638 11591 412694 11600
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 11591
rect 414308 480 414336 16546
rect 415412 1834 415440 79494
rect 419538 76936 419594 76945
rect 419538 76871 419594 76880
rect 417424 72480 417476 72486
rect 417424 72422 417476 72428
rect 417436 64394 417464 72422
rect 417424 64388 417476 64394
rect 417424 64330 417476 64336
rect 418160 49700 418212 49706
rect 418160 49642 418212 49648
rect 418172 46238 418200 49642
rect 418160 46232 418212 46238
rect 418160 46174 418212 46180
rect 416780 34332 416832 34338
rect 416780 34274 416832 34280
rect 415492 28688 415544 28694
rect 415492 28630 415544 28636
rect 415400 1828 415452 1834
rect 415400 1770 415452 1776
rect 415504 480 415532 28630
rect 416792 16574 416820 34274
rect 418160 21616 418212 21622
rect 418160 21558 418212 21564
rect 418172 16574 418200 21558
rect 419552 16574 419580 76871
rect 425060 69828 425112 69834
rect 425060 69770 425112 69776
rect 420184 68536 420236 68542
rect 420184 68478 420236 68484
rect 420196 36650 420224 68478
rect 422944 64388 422996 64394
rect 422944 64330 422996 64336
rect 422956 51882 422984 64330
rect 422944 51876 422996 51882
rect 422944 51818 422996 51824
rect 420184 36644 420236 36650
rect 420184 36586 420236 36592
rect 422300 34264 422352 34270
rect 422300 34206 422352 34212
rect 422312 16574 422340 34206
rect 423680 34196 423732 34202
rect 423680 34138 423732 34144
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 419552 16546 420224 16574
rect 422312 16546 422616 16574
rect 416688 1828 416740 1834
rect 416688 1770 416740 1776
rect 416700 480 416728 1770
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420196 480 420224 16546
rect 420920 14612 420972 14618
rect 420920 14554 420972 14560
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 14554
rect 422588 480 422616 16546
rect 423692 3398 423720 34138
rect 423772 31476 423824 31482
rect 423772 31418 423824 31424
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 423784 480 423812 31418
rect 425072 16574 425100 69770
rect 428464 51876 428516 51882
rect 428464 51818 428516 51824
rect 428476 36582 428504 51818
rect 429108 46232 429160 46238
rect 429108 46174 429160 46180
rect 429120 40730 429148 46174
rect 429108 40724 429160 40730
rect 429108 40666 429160 40672
rect 431960 39364 432012 39370
rect 431960 39306 432012 39312
rect 429844 36644 429896 36650
rect 429844 36586 429896 36592
rect 428464 36576 428516 36582
rect 428464 36518 428516 36524
rect 427820 34128 427872 34134
rect 427820 34070 427872 34076
rect 429198 34096 429254 34105
rect 426440 31408 426492 31414
rect 426440 31350 426492 31356
rect 426452 16574 426480 31350
rect 427832 16574 427860 34070
rect 429198 34031 429254 34040
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 427832 16546 428504 16574
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428476 480 428504 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 34031
rect 429856 32570 429884 36586
rect 429844 32564 429896 32570
rect 429844 32506 429896 32512
rect 430578 31376 430634 31385
rect 430578 31311 430634 31320
rect 430592 16574 430620 31311
rect 430592 16546 430896 16574
rect 430868 480 430896 16546
rect 431972 3398 432000 39306
rect 432050 33960 432106 33969
rect 432050 33895 432106 33904
rect 431960 3392 432012 3398
rect 431960 3334 432012 3340
rect 432064 480 432092 33895
rect 433352 16574 433380 80407
rect 462332 78985 462360 703520
rect 478524 700398 478552 703520
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494072 141438 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 494060 141432 494112 141438
rect 494060 141374 494112 141380
rect 526444 80164 526496 80170
rect 526444 80106 526496 80112
rect 462318 78976 462374 78985
rect 462318 78911 462374 78920
rect 454040 78464 454092 78470
rect 454040 78406 454092 78412
rect 451278 76800 451334 76809
rect 451278 76735 451334 76744
rect 446404 73840 446456 73846
rect 446404 73782 446456 73788
rect 445482 72448 445538 72457
rect 445482 72383 445538 72392
rect 445496 69290 445524 72383
rect 446416 69834 446444 73782
rect 446404 69828 446456 69834
rect 446404 69770 446456 69776
rect 445484 69284 445536 69290
rect 445484 69226 445536 69232
rect 447140 69284 447192 69290
rect 447140 69226 447192 69232
rect 439502 68232 439558 68241
rect 439502 68167 439558 68176
rect 437480 66904 437532 66910
rect 437480 66846 437532 66852
rect 434720 65544 434772 65550
rect 434720 65486 434772 65492
rect 434732 16574 434760 65486
rect 436100 17536 436152 17542
rect 436100 17478 436152 17484
rect 436112 16574 436140 17478
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 436112 16546 436784 16574
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 433260 480 433288 3334
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436756 480 436784 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 66846
rect 439516 62830 439544 68167
rect 447152 66230 447180 69226
rect 447140 66224 447192 66230
rect 447140 66166 447192 66172
rect 450636 66224 450688 66230
rect 450636 66166 450688 66172
rect 439504 62824 439556 62830
rect 439504 62766 439556 62772
rect 450648 60246 450676 66166
rect 450636 60240 450688 60246
rect 450636 60182 450688 60188
rect 440240 58744 440292 58750
rect 440240 58686 440292 58692
rect 439504 40724 439556 40730
rect 439504 40666 439556 40672
rect 438860 31340 438912 31346
rect 438860 31282 438912 31288
rect 438872 16574 438900 31282
rect 439516 26926 439544 40666
rect 439504 26920 439556 26926
rect 439504 26862 439556 26868
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 1834 440280 58686
rect 440332 49020 440384 49026
rect 440332 48962 440384 48968
rect 440240 1828 440292 1834
rect 440240 1770 440292 1776
rect 440344 480 440372 48962
rect 447140 43444 447192 43450
rect 447140 43386 447192 43392
rect 440884 32564 440936 32570
rect 440884 32506 440936 32512
rect 440896 24342 440924 32506
rect 446404 26920 446456 26926
rect 446404 26862 446456 26868
rect 440884 24336 440936 24342
rect 440884 24278 440936 24284
rect 443736 24336 443788 24342
rect 443736 24278 443788 24284
rect 443748 17950 443776 24278
rect 446416 22098 446444 26862
rect 446404 22092 446456 22098
rect 446404 22034 446456 22040
rect 443736 17944 443788 17950
rect 443736 17886 443788 17892
rect 444378 17776 444434 17785
rect 444378 17711 444434 17720
rect 441620 17468 441672 17474
rect 441620 17410 441672 17416
rect 441632 16574 441660 17410
rect 444392 16574 444420 17711
rect 445758 17640 445814 17649
rect 445758 17575 445814 17584
rect 441632 16546 442672 16574
rect 444392 16546 445064 16574
rect 441528 1828 441580 1834
rect 441528 1770 441580 1776
rect 441540 480 441568 1770
rect 442644 480 442672 16546
rect 443828 7608 443880 7614
rect 443828 7550 443880 7556
rect 443840 480 443868 7550
rect 445036 480 445064 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 17575
rect 447152 16574 447180 43386
rect 449900 28620 449952 28626
rect 449900 28562 449952 28568
rect 448888 22092 448940 22098
rect 448888 22034 448940 22040
rect 448900 18834 448928 22034
rect 448888 18828 448940 18834
rect 448888 18770 448940 18776
rect 449164 17944 449216 17950
rect 449164 17886 449216 17892
rect 448518 17504 448574 17513
rect 448518 17439 448574 17448
rect 448532 16574 448560 17439
rect 447152 16546 447456 16574
rect 448532 16546 448652 16574
rect 447428 480 447456 16546
rect 448624 480 448652 16546
rect 449176 14618 449204 17886
rect 449912 16574 449940 28562
rect 451292 16574 451320 76735
rect 452660 28552 452712 28558
rect 452660 28494 452712 28500
rect 449912 16546 450952 16574
rect 451292 16546 451688 16574
rect 449164 14612 449216 14618
rect 449164 14554 449216 14560
rect 449806 6216 449862 6225
rect 449806 6151 449862 6160
rect 449820 480 449848 6151
rect 450924 480 450952 16546
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 452672 6914 452700 28494
rect 452752 18828 452804 18834
rect 452752 18770 452804 18776
rect 452764 15638 452792 18770
rect 452752 15632 452804 15638
rect 452752 15574 452804 15580
rect 452672 6886 453344 6914
rect 453316 480 453344 6886
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 78406
rect 460940 78396 460992 78402
rect 460940 78338 460992 78344
rect 456064 71120 456116 71126
rect 456064 71062 456116 71068
rect 456076 43110 456104 71062
rect 460296 69828 460348 69834
rect 460296 69770 460348 69776
rect 460204 68468 460256 68474
rect 460204 68410 460256 68416
rect 458824 60240 458876 60246
rect 458824 60182 458876 60188
rect 458836 47598 458864 60182
rect 460216 57254 460244 68410
rect 460308 62898 460336 69770
rect 460296 62892 460348 62898
rect 460296 62834 460348 62840
rect 460204 57248 460256 57254
rect 460204 57190 460256 57196
rect 458824 47592 458876 47598
rect 458824 47534 458876 47540
rect 456064 43104 456116 43110
rect 456064 43046 456116 43052
rect 458548 43104 458600 43110
rect 458548 43046 458600 43052
rect 458560 36582 458588 43046
rect 454868 36576 454920 36582
rect 454868 36518 454920 36524
rect 458548 36576 458600 36582
rect 458548 36518 458600 36524
rect 454880 31414 454908 36518
rect 454868 31408 454920 31414
rect 454868 31350 454920 31356
rect 458824 31408 458876 31414
rect 458824 31350 458876 31356
rect 456892 28484 456944 28490
rect 456892 28426 456944 28432
rect 454592 14612 454644 14618
rect 454592 14554 454644 14560
rect 454604 7614 454632 14554
rect 455696 11824 455748 11830
rect 455696 11766 455748 11772
rect 454592 7608 454644 7614
rect 454592 7550 454644 7556
rect 455708 480 455736 11766
rect 456904 480 456932 28426
rect 458180 15632 458232 15638
rect 458180 15574 458232 15580
rect 458192 10402 458220 15574
rect 458836 12442 458864 31350
rect 459560 28416 459612 28422
rect 459560 28358 459612 28364
rect 459572 16574 459600 28358
rect 460952 16574 460980 78338
rect 467840 78328 467892 78334
rect 467840 78270 467892 78276
rect 467104 71052 467156 71058
rect 467104 70994 467156 71000
rect 464344 62892 464396 62898
rect 464344 62834 464396 62840
rect 463792 62824 463844 62830
rect 463792 62766 463844 62772
rect 463804 59430 463832 62766
rect 463792 59424 463844 59430
rect 463792 59366 463844 59372
rect 461308 47592 461360 47598
rect 461308 47534 461360 47540
rect 461320 40050 461348 47534
rect 461308 40044 461360 40050
rect 461308 39986 461360 39992
rect 463884 36576 463936 36582
rect 463884 36518 463936 36524
rect 463896 31346 463924 36518
rect 463884 31340 463936 31346
rect 463884 31282 463936 31288
rect 464356 26926 464384 62834
rect 464896 57248 464948 57254
rect 464896 57190 464948 57196
rect 464908 49706 464936 57190
rect 464896 49700 464948 49706
rect 464896 49642 464948 49648
rect 467116 33114 467144 70994
rect 467196 59424 467248 59430
rect 467196 59366 467248 59372
rect 467208 47598 467236 59366
rect 467196 47592 467248 47598
rect 467196 47534 467248 47540
rect 467104 33108 467156 33114
rect 467104 33050 467156 33056
rect 465078 31240 465134 31249
rect 465078 31175 465134 31184
rect 464344 26920 464396 26926
rect 464344 26862 464396 26868
rect 462320 17400 462372 17406
rect 462320 17342 462372 17348
rect 463698 17368 463754 17377
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 459192 14544 459244 14550
rect 459192 14486 459244 14492
rect 458824 12436 458876 12442
rect 458824 12378 458876 12384
rect 458180 10396 458232 10402
rect 458180 10338 458232 10344
rect 458088 3868 458140 3874
rect 458088 3810 458140 3816
rect 458100 480 458128 3810
rect 459204 480 459232 14486
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 461676 12436 461728 12442
rect 461676 12378 461728 12384
rect 461688 3874 461716 12378
rect 461676 3868 461728 3874
rect 461676 3810 461728 3816
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 17342
rect 463698 17303 463754 17312
rect 463712 16574 463740 17303
rect 463712 16546 464016 16574
rect 463988 480 464016 16546
rect 465092 6914 465120 31175
rect 466458 28384 466514 28393
rect 466458 28319 466514 28328
rect 465170 17232 465226 17241
rect 465170 17167 465226 17176
rect 465184 16574 465212 17167
rect 466472 16574 466500 28319
rect 467852 16574 467880 78270
rect 474740 78260 474792 78266
rect 474740 78202 474792 78208
rect 471244 49700 471296 49706
rect 471244 49642 471296 49648
rect 468484 40044 468536 40050
rect 468484 39986 468536 39992
rect 465184 16546 465672 16574
rect 466472 16546 467512 16574
rect 467852 16546 468248 16574
rect 465092 6886 465212 6914
rect 465184 480 465212 6886
rect 465644 490 465672 16546
rect 465724 10396 465776 10402
rect 465724 10338 465776 10344
rect 465736 3398 465764 10338
rect 465724 3392 465776 3398
rect 465724 3334 465776 3340
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465644 462 465856 490
rect 467484 480 467512 16546
rect 465828 354 465856 462
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468220 354 468248 16546
rect 468496 14550 468524 39986
rect 471256 34338 471284 49642
rect 471244 34332 471296 34338
rect 471244 34274 471296 34280
rect 472348 33108 472400 33114
rect 472348 33050 472400 33056
rect 472360 29714 472388 33050
rect 473360 31340 473412 31346
rect 473360 31282 473412 31288
rect 472348 29708 472400 29714
rect 472348 29650 472400 29656
rect 473372 16574 473400 31282
rect 474752 16574 474780 78202
rect 485780 75472 485832 75478
rect 485780 75414 485832 75420
rect 475382 69592 475438 69601
rect 475382 69527 475438 69536
rect 475396 62150 475424 69527
rect 475384 62144 475436 62150
rect 475384 62086 475436 62092
rect 479524 62144 479576 62150
rect 479524 62086 479576 62092
rect 478880 58676 478932 58682
rect 478880 58618 478932 58624
rect 476764 47592 476816 47598
rect 476764 47534 476816 47540
rect 476120 34332 476172 34338
rect 476120 34274 476172 34280
rect 476132 16574 476160 34274
rect 473372 16546 474136 16574
rect 474752 16546 475792 16574
rect 476132 16546 476528 16574
rect 468484 14544 468536 14550
rect 468484 14486 468536 14492
rect 473452 7608 473504 7614
rect 473452 7550 473504 7556
rect 471060 3868 471112 3874
rect 471060 3810 471112 3816
rect 469864 3392 469916 3398
rect 469864 3334 469916 3340
rect 469876 480 469904 3334
rect 471072 480 471100 3810
rect 472256 3800 472308 3806
rect 472256 3742 472308 3748
rect 472268 480 472296 3742
rect 473464 480 473492 7550
rect 468638 354 468750 480
rect 468220 326 468750 354
rect 468638 -960 468750 326
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 16546
rect 475764 480 475792 16546
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 16546
rect 476776 11830 476804 47534
rect 477500 29708 477552 29714
rect 477500 29650 477552 29656
rect 477512 16574 477540 29650
rect 477512 16546 478184 16574
rect 476764 11824 476816 11830
rect 476764 11766 476816 11772
rect 478156 480 478184 16546
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 478892 354 478920 58618
rect 479536 13802 479564 62086
rect 483018 31104 483074 31113
rect 483018 31039 483074 31048
rect 483032 16574 483060 31039
rect 485792 16574 485820 75414
rect 496820 75404 496872 75410
rect 496820 75346 496872 75352
rect 491300 60172 491352 60178
rect 491300 60114 491352 60120
rect 490012 29640 490064 29646
rect 490012 29582 490064 29588
rect 488540 20188 488592 20194
rect 488540 20130 488592 20136
rect 488552 16574 488580 20130
rect 483032 16546 484072 16574
rect 485792 16546 486464 16574
rect 488552 16546 488856 16574
rect 482284 14544 482336 14550
rect 482284 14486 482336 14492
rect 479524 13796 479576 13802
rect 479524 13738 479576 13744
rect 481732 13796 481784 13802
rect 481732 13738 481784 13744
rect 479524 11824 479576 11830
rect 479524 11766 479576 11772
rect 479536 5574 479564 11766
rect 479524 5568 479576 5574
rect 479524 5510 479576 5516
rect 480536 3732 480588 3738
rect 480536 3674 480588 3680
rect 480548 480 480576 3674
rect 481744 480 481772 13738
rect 482296 3194 482324 14486
rect 482836 5568 482888 5574
rect 482836 5510 482888 5516
rect 482284 3188 482336 3194
rect 482284 3130 482336 3136
rect 482848 480 482876 5510
rect 484044 480 484072 16546
rect 485228 3188 485280 3194
rect 485228 3130 485280 3136
rect 485240 480 485268 3130
rect 486436 480 486464 16546
rect 487620 3664 487672 3670
rect 487620 3606 487672 3612
rect 487632 480 487660 3606
rect 488828 480 488856 16546
rect 490024 6914 490052 29582
rect 491312 16574 491340 60114
rect 493324 26920 493376 26926
rect 493324 26862 493376 26868
rect 491312 16546 492352 16574
rect 489932 6886 490052 6914
rect 489932 480 489960 6886
rect 491116 3596 491168 3602
rect 491116 3538 491168 3544
rect 491128 480 491156 3538
rect 492324 480 492352 16546
rect 493336 13122 493364 26862
rect 495440 20120 495492 20126
rect 495440 20062 495492 20068
rect 493324 13116 493376 13122
rect 493324 13058 493376 13064
rect 493508 8968 493560 8974
rect 493508 8910 493560 8916
rect 493520 480 493548 8910
rect 494704 4888 494756 4894
rect 494704 4830 494756 4836
rect 494716 480 494744 4830
rect 479310 354 479422 480
rect 478892 326 479422 354
rect 479310 -960 479422 326
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495452 354 495480 20062
rect 496832 16574 496860 75346
rect 499580 75336 499632 75342
rect 499580 75278 499632 75284
rect 498200 68400 498252 68406
rect 498200 68342 498252 68348
rect 496832 16546 497136 16574
rect 497108 480 497136 16546
rect 498212 480 498240 68342
rect 498292 20052 498344 20058
rect 498292 19994 498344 20000
rect 498304 16574 498332 19994
rect 499592 16574 499620 75278
rect 514760 75268 514812 75274
rect 514760 75210 514812 75216
rect 500958 71224 501014 71233
rect 500958 71159 501014 71168
rect 500972 16574 501000 71159
rect 512000 69760 512052 69766
rect 512000 69702 512052 69708
rect 506480 25832 506532 25838
rect 506480 25774 506532 25780
rect 502338 21312 502394 21321
rect 502338 21247 502394 21256
rect 502352 16574 502380 21247
rect 498304 16546 498976 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 503720 10328 503772 10334
rect 503720 10270 503772 10276
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 10270
rect 506492 3534 506520 25774
rect 506572 21548 506624 21554
rect 506572 21490 506624 21496
rect 505376 3528 505428 3534
rect 505376 3470 505428 3476
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 505388 480 505416 3470
rect 506584 3346 506612 21490
rect 509240 21480 509292 21486
rect 509240 21422 509292 21428
rect 509252 16574 509280 21422
rect 509252 16546 509648 16574
rect 507860 13116 507912 13122
rect 507860 13058 507912 13064
rect 507872 8974 507900 13058
rect 507860 8968 507912 8974
rect 507860 8910 507912 8916
rect 507308 3528 507360 3534
rect 507308 3470 507360 3476
rect 506492 3318 506612 3346
rect 506492 480 506520 3318
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507320 354 507348 3470
rect 508872 3460 508924 3466
rect 508872 3402 508924 3408
rect 508884 480 508912 3402
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511264 11756 511316 11762
rect 511264 11698 511316 11704
rect 511276 480 511304 11698
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512012 354 512040 69702
rect 513380 21412 513432 21418
rect 513380 21354 513432 21360
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 21354
rect 514772 480 514800 75210
rect 518898 71088 518954 71097
rect 518898 71023 518954 71032
rect 514852 68332 514904 68338
rect 514852 68274 514904 68280
rect 514864 16574 514892 68274
rect 517518 24304 517574 24313
rect 517518 24239 517574 24248
rect 516138 22944 516194 22953
rect 516138 22879 516194 22888
rect 516152 16574 516180 22879
rect 517532 16574 517560 24239
rect 518912 16574 518940 71023
rect 521660 28348 521712 28354
rect 521660 28290 521712 28296
rect 520278 22808 520334 22817
rect 520278 22743 520334 22752
rect 514864 16546 515536 16574
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 518912 16546 519584 16574
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515508 354 515536 16546
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519556 480 519584 16546
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 22743
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 28290
rect 524420 28280 524472 28286
rect 524420 28222 524472 28228
rect 523040 17332 523092 17338
rect 523040 17274 523092 17280
rect 523052 16574 523080 17274
rect 524432 16574 524460 28222
rect 526456 20670 526484 80106
rect 527192 79354 527220 703520
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 558932 140078 558960 702406
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580538 670712 580594 670721
rect 580538 670647 580594 670656
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 580262 591016 580318 591025
rect 580262 590951 580318 590960
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 576910 579660 577623
rect 579620 576904 579672 576910
rect 579620 576846 579672 576852
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 579802 524512 579858 524521
rect 579802 524447 579804 524456
rect 579856 524447 579858 524456
rect 579804 524418 579856 524424
rect 579986 511320 580042 511329
rect 579986 511255 580042 511264
rect 580000 510678 580028 511255
rect 579988 510672 580040 510678
rect 579988 510614 580040 510620
rect 579618 471472 579674 471481
rect 579618 471407 579674 471416
rect 579632 470626 579660 471407
rect 579620 470620 579672 470626
rect 579620 470562 579672 470568
rect 579618 458144 579674 458153
rect 579618 458079 579674 458088
rect 579632 456822 579660 458079
rect 579620 456816 579672 456822
rect 579620 456758 579672 456764
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579724 418198 579752 418231
rect 579712 418192 579764 418198
rect 579712 418134 579764 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244322 580212 245511
rect 580172 244316 580224 244322
rect 580172 244258 580224 244264
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 579986 219056 580042 219065
rect 579986 218991 580042 219000
rect 580000 218074 580028 218991
rect 579988 218068 580040 218074
rect 579988 218010 580040 218016
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 558920 140072 558972 140078
rect 558920 140014 558972 140020
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580078 112840 580134 112849
rect 580078 112775 580134 112784
rect 580092 111858 580120 112775
rect 580080 111852 580132 111858
rect 580080 111794 580132 111800
rect 579986 99512 580042 99521
rect 579986 99447 580042 99456
rect 580000 94518 580028 99447
rect 580184 94586 580212 139295
rect 580172 94580 580224 94586
rect 580172 94522 580224 94528
rect 579988 94512 580040 94518
rect 579988 94454 580040 94460
rect 580172 86420 580224 86426
rect 580172 86362 580224 86368
rect 527180 79348 527232 79354
rect 527180 79290 527232 79296
rect 557540 78192 557592 78198
rect 557540 78134 557592 78140
rect 535458 76664 535514 76673
rect 535458 76599 535514 76608
rect 529940 60104 529992 60110
rect 529940 60046 529992 60052
rect 528560 25764 528612 25770
rect 528560 25706 528612 25712
rect 526444 20664 526496 20670
rect 526444 20606 526496 20612
rect 527180 17264 527232 17270
rect 527180 17206 527232 17212
rect 527192 16574 527220 17206
rect 523052 16546 523816 16574
rect 524432 16546 525472 16574
rect 527192 16546 527864 16574
rect 523038 3496 523094 3505
rect 523038 3431 523094 3440
rect 523052 480 523080 3431
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525444 480 525472 16546
rect 526628 8968 526680 8974
rect 526628 8910 526680 8916
rect 526640 480 526668 8910
rect 527836 480 527864 16546
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 25706
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 60046
rect 531318 28248 531374 28257
rect 531318 28183 531374 28192
rect 531332 3534 531360 28183
rect 531412 19984 531464 19990
rect 531412 19926 531464 19932
rect 534078 19952 534134 19961
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531424 3346 531452 19926
rect 534078 19887 534134 19896
rect 534092 16574 534120 19887
rect 535472 16574 535500 76599
rect 549258 76528 549314 76537
rect 549258 76463 549314 76472
rect 547878 75304 547934 75313
rect 547878 75239 547934 75248
rect 543740 75200 543792 75206
rect 543740 75142 543792 75148
rect 539600 69692 539652 69698
rect 539600 69634 539652 69640
rect 536838 61568 536894 61577
rect 536838 61503 536894 61512
rect 536852 16574 536880 61503
rect 538218 22672 538274 22681
rect 538218 22607 538274 22616
rect 534092 16546 534488 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 533712 4820 533764 4826
rect 533712 4762 533764 4768
rect 532148 3528 532200 3534
rect 532148 3470 532200 3476
rect 531332 3318 531452 3346
rect 531332 480 531360 3318
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3470
rect 533724 480 533752 4762
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 22607
rect 539612 3534 539640 69634
rect 539692 34060 539744 34066
rect 539692 34002 539744 34008
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 34002
rect 542360 33992 542412 33998
rect 542360 33934 542412 33940
rect 540980 31272 541032 31278
rect 540980 31214 541032 31220
rect 540992 16574 541020 31214
rect 542372 16574 542400 33934
rect 543752 16574 543780 75142
rect 546500 33924 546552 33930
rect 546500 33866 546552 33872
rect 545120 31204 545172 31210
rect 545120 31146 545172 31152
rect 545132 16574 545160 31146
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 33866
rect 547892 480 547920 75239
rect 547972 31136 548024 31142
rect 547972 31078 548024 31084
rect 547984 16574 548012 31078
rect 549272 16574 549300 76463
rect 552020 33856 552072 33862
rect 552020 33798 552072 33804
rect 556158 33824 556214 33833
rect 550640 31068 550692 31074
rect 550640 31010 550692 31016
rect 550652 16574 550680 31010
rect 552032 16574 552060 33798
rect 553400 33788 553452 33794
rect 556158 33759 556214 33768
rect 553400 33730 553452 33736
rect 553412 16574 553440 33730
rect 554778 30968 554834 30977
rect 554778 30903 554834 30912
rect 547984 16546 548656 16574
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 553412 16546 553808 16574
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 550284 480 550312 16546
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 30903
rect 556172 480 556200 33759
rect 556252 32496 556304 32502
rect 556252 32438 556304 32444
rect 556264 16574 556292 32438
rect 557552 16574 557580 78134
rect 574100 78124 574152 78130
rect 574100 78066 574152 78072
rect 571338 75168 571394 75177
rect 571338 75103 571394 75112
rect 568580 64184 568632 64190
rect 568580 64126 568632 64132
rect 564440 60036 564492 60042
rect 564440 59978 564492 59984
rect 558920 25696 558972 25702
rect 558920 25638 558972 25644
rect 558932 16574 558960 25638
rect 563060 25628 563112 25634
rect 563060 25570 563112 25576
rect 560300 18624 560352 18630
rect 560300 18566 560352 18572
rect 560312 16574 560340 18566
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562046 3360 562102 3369
rect 562046 3295 562102 3304
rect 562060 480 562088 3295
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 25570
rect 564452 3534 564480 59978
rect 564532 32428 564584 32434
rect 564532 32370 564584 32376
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 32370
rect 565820 25560 565872 25566
rect 565820 25502 565872 25508
rect 565832 16574 565860 25502
rect 568592 16574 568620 64126
rect 569958 24168 570014 24177
rect 569958 24103 570014 24112
rect 569972 16574 570000 24103
rect 565832 16546 566872 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566844 480 566872 16546
rect 567568 14476 567620 14482
rect 567568 14418 567620 14424
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 14418
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571352 354 571380 75103
rect 572718 62928 572774 62937
rect 572718 62863 572774 62872
rect 572732 480 572760 62863
rect 574112 16574 574140 78066
rect 580184 77926 580212 86362
rect 580276 80782 580304 590951
rect 580354 537840 580410 537849
rect 580354 537775 580410 537784
rect 580264 80776 580316 80782
rect 580264 80718 580316 80724
rect 580368 80714 580396 537775
rect 580552 485110 580580 670647
rect 580540 485104 580592 485110
rect 580540 485046 580592 485052
rect 580446 484664 580502 484673
rect 580446 484599 580502 484608
rect 580356 80708 580408 80714
rect 580356 80650 580408 80656
rect 580460 80102 580488 484599
rect 580538 431624 580594 431633
rect 580538 431559 580594 431568
rect 580448 80096 580500 80102
rect 580448 80038 580500 80044
rect 580552 78849 580580 431559
rect 580630 378448 580686 378457
rect 580630 378383 580686 378392
rect 580538 78840 580594 78849
rect 580538 78775 580594 78784
rect 580644 78606 580672 378383
rect 580722 325272 580778 325281
rect 580722 325207 580778 325216
rect 580736 78713 580764 325207
rect 580814 272232 580870 272241
rect 580814 272167 580870 272176
rect 580828 86426 580856 272167
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 580816 86420 580868 86426
rect 580816 86362 580868 86368
rect 580814 86184 580870 86193
rect 580814 86119 580870 86128
rect 580828 80617 580856 86119
rect 580814 80608 580870 80617
rect 580814 80543 580870 80552
rect 580722 78704 580778 78713
rect 580722 78639 580778 78648
rect 580632 78600 580684 78606
rect 580632 78542 580684 78548
rect 580172 77920 580224 77926
rect 580172 77862 580224 77868
rect 580920 75886 580948 125967
rect 581000 78056 581052 78062
rect 581000 77998 581052 78004
rect 580908 75880 580960 75886
rect 580908 75822 580960 75828
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 575478 61432 575534 61441
rect 575478 61367 575534 61376
rect 575492 16574 575520 61367
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 576858 46200 576914 46209
rect 576858 46135 576914 46144
rect 576872 16574 576900 46135
rect 580264 44872 580316 44878
rect 580264 44814 580316 44820
rect 580276 33153 580304 44814
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 580264 22772 580316 22778
rect 580264 22714 580316 22720
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 574112 16546 575152 16574
rect 575492 16546 575888 16574
rect 576872 16546 576992 16574
rect 573916 6248 573968 6254
rect 573916 6190 573968 6196
rect 573928 480 573956 6190
rect 575124 480 575152 16546
rect 571494 354 571606 480
rect 571352 326 571606 354
rect 571494 -960 571606 326
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 575860 354 575888 16546
rect 576278 354 576390 480
rect 575860 326 576390 354
rect 576964 354 576992 16546
rect 580276 6633 580304 22714
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 578608 6180 578660 6186
rect 578608 6122 578660 6128
rect 578620 480 578648 6122
rect 581012 480 581040 77998
rect 582380 77988 582432 77994
rect 582380 77930 582432 77936
rect 581090 62792 581146 62801
rect 581090 62727 581146 62736
rect 581104 16574 581132 62727
rect 582392 16574 582420 77930
rect 581104 16546 581776 16574
rect 582392 16546 583432 16574
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 576278 -960 576390 326
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583404 480 583432 16546
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3422 606056 3478 606112
rect 3330 579944 3386 580000
rect 3330 553832 3386 553888
rect 3330 527876 3386 527912
rect 3330 527856 3332 527876
rect 3332 527856 3384 527876
rect 3384 527856 3386 527876
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3054 462576 3110 462632
rect 2962 449520 3018 449576
rect 3330 423544 3386 423600
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 3330 345344 3386 345400
rect 3146 319232 3202 319288
rect 3330 306176 3386 306232
rect 3238 267144 3294 267200
rect 2870 254088 2926 254144
rect 3330 214920 3386 214976
rect 3330 201864 3386 201920
rect 3330 188808 3386 188864
rect 3330 162868 3332 162888
rect 3332 162868 3384 162888
rect 3384 162868 3386 162888
rect 3330 162832 3386 162868
rect 3330 110608 3386 110664
rect 3330 84632 3386 84688
rect 3606 619112 3662 619168
rect 3514 149776 3570 149832
rect 3790 566888 3846 566944
rect 3698 501744 3754 501800
rect 3514 136720 3570 136776
rect 3514 97552 3570 97608
rect 3882 475632 3938 475688
rect 3882 358400 3938 358456
rect 3974 293120 4030 293176
rect 4066 241032 4122 241088
rect 3422 79192 3478 79248
rect 6918 79600 6974 79656
rect 4066 78512 4122 78568
rect 6918 75112 6974 75168
rect 3422 71612 3424 71632
rect 3424 71612 3476 71632
rect 3476 71612 3478 71632
rect 3422 71576 3478 71612
rect 3422 58520 3478 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 32408 3478 32464
rect 2962 19352 3018 19408
rect 3422 6432 3478 6488
rect 8298 72392 8354 72448
rect 71778 79464 71834 79520
rect 117318 137536 117374 137592
rect 117318 136040 117374 136096
rect 117318 134544 117374 134600
rect 117410 133048 117466 133104
rect 117318 131552 117374 131608
rect 117318 130056 117374 130112
rect 117318 128560 117374 128616
rect 117318 127064 117374 127120
rect 117318 125568 117374 125624
rect 117318 124108 117320 124128
rect 117320 124108 117372 124128
rect 117372 124108 117374 124128
rect 117318 124072 117374 124108
rect 117318 122576 117374 122632
rect 117318 121080 117374 121136
rect 117318 119584 117374 119640
rect 117318 118088 117374 118144
rect 117318 116592 117374 116648
rect 117318 115096 117374 115152
rect 118054 113600 118110 113656
rect 118238 92656 118294 92712
rect 118146 91160 118202 91216
rect 118974 110608 119030 110664
rect 119066 109112 119122 109168
rect 119250 112104 119306 112160
rect 119158 107616 119214 107672
rect 118882 106120 118938 106176
rect 118790 104624 118846 104680
rect 118698 103128 118754 103184
rect 118606 95648 118662 95704
rect 118514 94152 118570 94208
rect 118422 89664 118478 89720
rect 118330 88168 118386 88224
rect 118514 86672 118570 86728
rect 118422 83680 118478 83736
rect 116582 79328 116638 79384
rect 27618 72528 27674 72584
rect 11150 35128 11206 35184
rect 26514 6296 26570 6352
rect 25318 6160 25374 6216
rect 46938 75248 46994 75304
rect 45466 8880 45522 8936
rect 44270 7520 44326 7576
rect 48962 7656 49018 7712
rect 64878 73752 64934 73808
rect 60738 22616 60794 22672
rect 64326 7928 64382 7984
rect 63222 7792 63278 7848
rect 95882 77832 95938 77888
rect 80058 75384 80114 75440
rect 78126 10240 78182 10296
rect 88890 6432 88946 6488
rect 95790 10376 95846 10432
rect 97998 72664 98054 72720
rect 115938 76472 115994 76528
rect 101034 3304 101090 3360
rect 114006 11600 114062 11656
rect 118606 85176 118662 85232
rect 118606 80552 118662 80608
rect 120722 102040 120778 102096
rect 120814 100680 120870 100736
rect 120906 98640 120962 98696
rect 120998 97144 121054 97200
rect 120722 81640 120778 81696
rect 119342 78376 119398 78432
rect 119894 9016 119950 9072
rect 124862 77968 124918 78024
rect 126886 75112 126942 75168
rect 129646 77696 129702 77752
rect 130106 79872 130162 79928
rect 131072 79906 131128 79962
rect 131440 79906 131496 79962
rect 131808 79906 131864 79962
rect 132176 79906 132232 79962
rect 132360 79906 132416 79962
rect 130750 72528 130806 72584
rect 131762 79736 131818 79792
rect 131026 77152 131082 77208
rect 131394 78104 131450 78160
rect 131118 73208 131174 73264
rect 132222 79736 132278 79792
rect 132728 79872 132784 79928
rect 132912 79906 132968 79962
rect 132682 79736 132738 79792
rect 133280 79906 133336 79962
rect 133464 79872 133520 79928
rect 133648 79906 133704 79962
rect 133234 79736 133290 79792
rect 133418 79736 133474 79792
rect 132406 75248 132462 75304
rect 132866 78104 132922 78160
rect 132590 75792 132646 75848
rect 133326 77968 133382 78024
rect 133602 79736 133658 79792
rect 134016 79906 134072 79962
rect 134062 79736 134118 79792
rect 133970 78648 134026 78704
rect 134384 79736 134440 79792
rect 135028 79872 135084 79928
rect 135258 79736 135314 79792
rect 135488 79872 135544 79928
rect 135074 78648 135130 78704
rect 135672 79736 135728 79792
rect 135534 77288 135590 77344
rect 135902 79056 135958 79112
rect 136500 79872 136556 79928
rect 136638 79736 136694 79792
rect 136270 78784 136326 78840
rect 136178 78648 136234 78704
rect 136730 78648 136786 78704
rect 137052 79872 137108 79928
rect 137144 79736 137200 79792
rect 136730 77832 136786 77888
rect 137742 78784 137798 78840
rect 137742 78648 137798 78704
rect 138340 79906 138396 79962
rect 138294 79736 138350 79792
rect 138524 79872 138580 79928
rect 138202 78920 138258 78976
rect 138110 78648 138166 78704
rect 138386 78784 138442 78840
rect 138984 79872 139040 79928
rect 138938 79736 138994 79792
rect 139628 79906 139684 79962
rect 139904 79872 139960 79928
rect 140272 79906 140328 79962
rect 140732 79872 140788 79928
rect 140134 79736 140190 79792
rect 139490 78648 139546 78704
rect 140594 79736 140650 79792
rect 141192 79770 141248 79826
rect 140870 77580 140926 77616
rect 140870 77560 140872 77580
rect 140872 77560 140924 77580
rect 140924 77560 140926 77580
rect 141652 79872 141708 79928
rect 142664 79872 142720 79928
rect 141238 78648 141294 78704
rect 142066 76608 142122 76664
rect 142342 76608 142398 76664
rect 143492 79872 143548 79928
rect 143676 79906 143732 79962
rect 143446 79736 143502 79792
rect 143354 77424 143410 77480
rect 143262 77288 143318 77344
rect 144228 79872 144284 79928
rect 144688 79872 144744 79928
rect 144826 79772 144828 79792
rect 144828 79772 144880 79792
rect 144880 79772 144882 79792
rect 144090 77560 144146 77616
rect 144550 77424 144606 77480
rect 144550 76608 144606 76664
rect 144826 79736 144882 79772
rect 144918 77424 144974 77480
rect 145884 79872 145940 79928
rect 145654 77424 145710 77480
rect 146206 77424 146262 77480
rect 146528 79736 146584 79792
rect 147080 79872 147136 79928
rect 147448 79906 147504 79962
rect 146574 77288 146630 77344
rect 146666 76608 146722 76664
rect 148460 79906 148516 79962
rect 148644 79906 148700 79962
rect 148828 79872 148884 79928
rect 149104 79906 149160 79962
rect 147494 77424 147550 77480
rect 147402 77288 147458 77344
rect 149564 79906 149620 79962
rect 149748 79872 149804 79928
rect 148046 76608 148102 76664
rect 149058 79736 149114 79792
rect 148782 76064 148838 76120
rect 148874 75928 148930 75984
rect 148322 3576 148378 3632
rect 149242 79056 149298 79112
rect 149426 76744 149482 76800
rect 149426 76064 149482 76120
rect 150300 79906 150356 79962
rect 150760 79906 150816 79962
rect 149702 75928 149758 75984
rect 150944 79906 151000 79962
rect 151680 79906 151736 79962
rect 150070 76608 150126 76664
rect 149978 75928 150034 75984
rect 150254 74024 150310 74080
rect 150990 78240 151046 78296
rect 150070 3712 150126 3768
rect 150714 75928 150770 75984
rect 151266 78104 151322 78160
rect 152324 79906 152380 79962
rect 152692 79872 152748 79928
rect 152876 79906 152932 79962
rect 153428 79906 153484 79962
rect 153704 79872 153760 79928
rect 151634 75928 151690 75984
rect 152186 77152 152242 77208
rect 152186 75928 152242 75984
rect 153106 76064 153162 76120
rect 152830 75928 152886 75984
rect 154440 79906 154496 79962
rect 154900 79872 154956 79928
rect 155360 79906 155416 79962
rect 155544 79906 155600 79962
rect 153566 75928 153622 75984
rect 153750 77016 153806 77072
rect 154394 77696 154450 77752
rect 154302 77016 154358 77072
rect 154486 75928 154542 75984
rect 155314 79736 155370 79792
rect 155820 79906 155876 79962
rect 156464 79906 156520 79962
rect 156740 79872 156796 79928
rect 156648 79736 156704 79792
rect 155682 75656 155738 75712
rect 156694 78920 156750 78976
rect 157752 79906 157808 79962
rect 157936 79906 157992 79962
rect 158488 79872 158544 79928
rect 157016 79736 157072 79792
rect 158580 79772 158582 79792
rect 158582 79772 158634 79792
rect 158634 79772 158636 79792
rect 156786 75520 156842 75576
rect 156970 75928 157026 75984
rect 156878 75384 156934 75440
rect 157154 76064 157210 76120
rect 157430 79056 157486 79112
rect 157706 79600 157762 79656
rect 157614 74296 157670 74352
rect 157246 73888 157302 73944
rect 157614 73772 157670 73808
rect 157614 73752 157616 73772
rect 157616 73752 157668 73772
rect 157668 73752 157670 73772
rect 158350 79600 158406 79656
rect 158580 79736 158636 79772
rect 159316 79872 159372 79928
rect 158626 78920 158682 78976
rect 160512 79906 160568 79962
rect 158442 76880 158498 76936
rect 158258 76200 158314 76256
rect 158626 73752 158682 73808
rect 159270 79600 159326 79656
rect 159638 79600 159694 79656
rect 160972 79872 161028 79928
rect 161340 79906 161396 79962
rect 160098 76880 160154 76936
rect 160006 74840 160062 74896
rect 150530 3576 150586 3632
rect 161110 79736 161166 79792
rect 161616 79872 161672 79928
rect 161984 79906 162040 79962
rect 162352 79906 162408 79962
rect 161202 79600 161258 79656
rect 161110 78784 161166 78840
rect 161294 77288 161350 77344
rect 161570 78784 161626 78840
rect 161938 78784 161994 78840
rect 161846 78648 161902 78704
rect 162444 79736 162500 79792
rect 162306 78920 162362 78976
rect 162720 79906 162776 79962
rect 163180 79872 163236 79928
rect 162490 78648 162546 78704
rect 162858 79056 162914 79112
rect 163640 79906 163696 79962
rect 164100 79872 164156 79928
rect 164376 79906 164432 79962
rect 163594 79636 163596 79656
rect 163596 79636 163648 79656
rect 163648 79636 163650 79656
rect 163594 79600 163650 79636
rect 163502 79056 163558 79112
rect 163318 78648 163374 78704
rect 163594 76880 163650 76936
rect 164054 78920 164110 78976
rect 163962 78648 164018 78704
rect 164146 78784 164202 78840
rect 164744 79872 164800 79928
rect 165204 79872 165260 79928
rect 164514 79600 164570 79656
rect 164422 78920 164478 78976
rect 162950 18672 163006 18728
rect 162490 4936 162546 4992
rect 165480 79872 165536 79928
rect 165250 78648 165306 78704
rect 165618 79056 165674 79112
rect 165526 78648 165582 78704
rect 165434 77968 165490 78024
rect 166584 79872 166640 79928
rect 167044 79872 167100 79928
rect 167504 79872 167560 79928
rect 167688 79906 167744 79962
rect 166630 79600 166686 79656
rect 166446 78784 166502 78840
rect 166722 78784 166778 78840
rect 166906 78648 166962 78704
rect 166814 78240 166870 78296
rect 166078 4800 166134 4856
rect 164882 3440 164938 3496
rect 167366 79600 167422 79656
rect 167642 79600 167698 79656
rect 167550 78104 167606 78160
rect 168332 79906 168388 79962
rect 168102 79600 168158 79656
rect 168102 79056 168158 79112
rect 168286 78920 168342 78976
rect 168194 78648 168250 78704
rect 168010 77560 168066 77616
rect 168700 79872 168756 79928
rect 168746 79736 168802 79792
rect 168562 79464 168618 79520
rect 168562 79076 168618 79112
rect 168562 79056 168564 79076
rect 168564 79056 168616 79076
rect 168616 79056 168618 79076
rect 168654 75928 168710 75984
rect 169160 79872 169216 79928
rect 169712 79872 169768 79928
rect 170080 79906 170136 79962
rect 170356 79906 170412 79962
rect 169666 78648 169722 78704
rect 168378 3304 168434 3360
rect 170402 79736 170458 79792
rect 170494 79464 170550 79520
rect 170402 77152 170458 77208
rect 170218 75928 170274 75984
rect 170678 77832 170734 77888
rect 171000 79872 171056 79928
rect 171276 79872 171332 79928
rect 171736 79906 171792 79962
rect 172012 79772 172014 79792
rect 172014 79772 172066 79792
rect 172066 79772 172068 79792
rect 171046 78648 171102 78704
rect 170954 78376 171010 78432
rect 170954 77696 171010 77752
rect 170862 75928 170918 75984
rect 172012 79736 172068 79772
rect 172518 79736 172574 79792
rect 171782 75928 171838 75984
rect 172426 79464 172482 79520
rect 172150 78648 172206 78704
rect 172150 78512 172206 78568
rect 172334 78376 172390 78432
rect 172242 76336 172298 76392
rect 171782 28192 171838 28248
rect 173392 79872 173448 79928
rect 173760 79906 173816 79962
rect 174128 79906 174184 79962
rect 174680 79872 174736 79928
rect 174956 79872 175012 79928
rect 175232 79906 175288 79962
rect 175416 79906 175472 79962
rect 173346 79464 173402 79520
rect 173714 77288 173770 77344
rect 174772 79772 174774 79792
rect 174774 79772 174826 79792
rect 174826 79772 174828 79792
rect 174174 78512 174230 78568
rect 174266 78376 174322 78432
rect 174174 77832 174230 77888
rect 174772 79736 174828 79772
rect 174910 79736 174966 79792
rect 174634 77832 174690 77888
rect 175002 76472 175058 76528
rect 175186 79056 175242 79112
rect 175186 78648 175242 78704
rect 175094 75248 175150 75304
rect 175784 79906 175840 79962
rect 175554 78376 175610 78432
rect 176428 79872 176484 79928
rect 177164 79872 177220 79928
rect 176014 78648 176070 78704
rect 175462 75928 175518 75984
rect 175370 75248 175426 75304
rect 177118 79736 177174 79792
rect 176658 78784 176714 78840
rect 176566 78648 176622 78704
rect 176290 76744 176346 76800
rect 176474 77696 176530 77752
rect 176474 77424 176530 77480
rect 176474 73480 176530 73536
rect 176934 78784 176990 78840
rect 177210 79328 177266 79384
rect 177118 79056 177174 79112
rect 177026 78240 177082 78296
rect 177992 79872 178048 79928
rect 177946 79736 178002 79792
rect 178544 79872 178600 79928
rect 178038 79600 178094 79656
rect 177670 79464 177726 79520
rect 177486 79056 177542 79112
rect 178222 79192 178278 79248
rect 177118 78104 177174 78160
rect 176842 77288 176898 77344
rect 177578 77696 177634 77752
rect 177394 75792 177450 75848
rect 178406 79192 178462 79248
rect 178498 78920 178554 78976
rect 179096 79906 179152 79962
rect 178314 78104 178370 78160
rect 178038 77968 178094 78024
rect 179050 77424 179106 77480
rect 178958 74840 179014 74896
rect 178866 74160 178922 74216
rect 179694 78376 179750 78432
rect 179878 78512 179934 78568
rect 180614 79736 180670 79792
rect 180522 78920 180578 78976
rect 188986 78240 189042 78296
rect 189078 77288 189134 77344
rect 181442 76608 181498 76664
rect 181442 76336 181498 76392
rect 179418 74976 179474 75032
rect 179418 68448 179474 68504
rect 182178 66816 182234 66872
rect 183558 57160 183614 57216
rect 189354 120672 189410 120728
rect 189354 116592 189410 116648
rect 189446 113872 189502 113928
rect 189630 130464 189686 130520
rect 189630 126112 189686 126168
rect 189722 119312 189778 119368
rect 189538 112512 189594 112568
rect 189354 82320 189410 82376
rect 189354 77560 189410 77616
rect 190734 129648 190790 129704
rect 190642 124208 190698 124264
rect 190550 117408 190606 117464
rect 190826 114688 190882 114744
rect 191930 128288 191986 128344
rect 191194 126928 191250 126984
rect 192022 122848 192078 122904
rect 191102 121488 191158 121544
rect 191010 110608 191066 110664
rect 190918 109248 190974 109304
rect 191930 107888 191986 107944
rect 191930 106528 191986 106584
rect 191930 105168 191986 105224
rect 191930 101124 191932 101144
rect 191932 101124 191984 101144
rect 191984 101124 191986 101144
rect 191930 101088 191986 101124
rect 192390 99728 192446 99784
rect 192114 98368 192170 98424
rect 192206 97008 192262 97064
rect 191930 95648 191986 95704
rect 192574 92928 192630 92984
rect 192574 82048 192630 82104
rect 193126 103808 193182 103864
rect 193126 102484 193128 102504
rect 193128 102484 193180 102504
rect 193180 102484 193182 102504
rect 193126 102448 193182 102484
rect 193126 94288 193182 94344
rect 193126 91568 193182 91624
rect 193126 90208 193182 90264
rect 193126 88848 193182 88904
rect 192942 87488 192998 87544
rect 193034 86128 193090 86184
rect 193126 84768 193182 84824
rect 193126 83408 193182 83464
rect 193126 80688 193182 80744
rect 331218 79464 331274 79520
rect 433338 80416 433394 80472
rect 397458 79056 397514 79112
rect 200118 63008 200174 63064
rect 201590 25472 201646 25528
rect 216678 34176 216734 34232
rect 215298 23296 215354 23352
rect 218150 6024 218206 6080
rect 303618 77016 303674 77072
rect 251178 74024 251234 74080
rect 241518 20440 241574 20496
rect 234618 18536 234674 18592
rect 232226 3984 232282 4040
rect 236550 10376 236606 10432
rect 235814 3848 235870 3904
rect 242990 3712 243046 3768
rect 249982 6840 250038 6896
rect 251270 12008 251326 12064
rect 253478 6704 253534 6760
rect 261574 71712 261630 71768
rect 266358 20304 266414 20360
rect 272890 75656 272946 75712
rect 264150 3576 264206 3632
rect 272430 11872 272486 11928
rect 271234 6568 271290 6624
rect 280894 71576 280950 71632
rect 289174 72528 289230 72584
rect 295338 73888 295394 73944
rect 284298 23160 284354 23216
rect 287058 23024 287114 23080
rect 286598 14456 286654 14512
rect 285402 6432 285458 6488
rect 288990 6296 289046 6352
rect 292578 28464 292634 28520
rect 303250 68312 303306 68368
rect 305642 75520 305698 75576
rect 310242 75384 310298 75440
rect 318154 73752 318210 73808
rect 310426 71440 310482 71496
rect 303158 9152 303214 9208
rect 306746 9016 306802 9072
rect 307942 8880 307998 8936
rect 396078 71304 396134 71360
rect 394698 48864 394754 48920
rect 392582 10240 392638 10296
rect 409878 20168 409934 20224
rect 414018 20032 414074 20088
rect 409142 11736 409198 11792
rect 412638 11600 412694 11656
rect 419538 76880 419594 76936
rect 429198 34040 429254 34096
rect 430578 31320 430634 31376
rect 432050 33904 432106 33960
rect 462318 78920 462374 78976
rect 451278 76744 451334 76800
rect 445482 72392 445538 72448
rect 439502 68176 439558 68232
rect 444378 17720 444434 17776
rect 445758 17584 445814 17640
rect 448518 17448 448574 17504
rect 449806 6160 449862 6216
rect 465078 31184 465134 31240
rect 463698 17312 463754 17368
rect 466458 28328 466514 28384
rect 465170 17176 465226 17232
rect 475382 69536 475438 69592
rect 483018 31048 483074 31104
rect 500958 71168 501014 71224
rect 502338 21256 502394 21312
rect 518898 71032 518954 71088
rect 517518 24248 517574 24304
rect 516138 22888 516194 22944
rect 520278 22752 520334 22808
rect 580170 683848 580226 683904
rect 580538 670656 580594 670712
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 580262 590960 580318 591016
rect 579618 577632 579674 577688
rect 580170 564304 580226 564360
rect 579802 524476 579858 524512
rect 579802 524456 579804 524476
rect 579804 524456 579856 524476
rect 579856 524456 579858 524476
rect 579986 511264 580042 511320
rect 579618 471416 579674 471472
rect 579618 458088 579674 458144
rect 579710 418240 579766 418296
rect 580170 404912 580226 404968
rect 580170 365064 580226 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 258848 580226 258904
rect 580170 245520 580226 245576
rect 579802 232328 579858 232384
rect 579986 219000 580042 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 579986 152632 580042 152688
rect 580170 139304 580226 139360
rect 580078 112784 580134 112840
rect 579986 99456 580042 99512
rect 535458 76608 535514 76664
rect 523038 3440 523094 3496
rect 531318 28192 531374 28248
rect 534078 19896 534134 19952
rect 549258 76472 549314 76528
rect 547878 75248 547934 75304
rect 536838 61512 536894 61568
rect 538218 22616 538274 22672
rect 556158 33768 556214 33824
rect 554778 30912 554834 30968
rect 571338 75112 571394 75168
rect 562046 3304 562102 3360
rect 569958 24112 570014 24168
rect 572718 62872 572774 62928
rect 580354 537784 580410 537840
rect 580446 484608 580502 484664
rect 580538 431568 580594 431624
rect 580630 378392 580686 378448
rect 580538 78784 580594 78840
rect 580722 325216 580778 325272
rect 580814 272176 580870 272232
rect 580906 125976 580962 126032
rect 580814 86128 580870 86184
rect 580814 80552 580870 80608
rect 580722 78648 580778 78704
rect 580170 72936 580226 72992
rect 575478 61376 575534 61432
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 576858 46144 576914 46200
rect 580262 33088 580318 33144
rect 579986 19760 580042 19816
rect 580262 6568 580318 6624
rect 581090 62736 581146 62792
<< metal3 >>
rect -960 697220 480 697460
rect 580206 697172 580212 697236
rect 580276 697234 580282 697236
rect 583520 697234 584960 697324
rect 580276 697174 584960 697234
rect 580276 697172 580282 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580533 670714 580599 670717
rect 583520 670714 584960 670804
rect 580533 670712 584960 670714
rect 580533 670656 580538 670712
rect 580594 670656 584960 670712
rect 580533 670654 584960 670656
rect 580533 670651 580599 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580390 643996 580396 644060
rect 580460 644058 580466 644060
rect 583520 644058 584960 644148
rect 580460 643998 584960 644058
rect 580460 643996 580466 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3601 619170 3667 619173
rect -960 619168 3667 619170
rect -960 619112 3606 619168
rect 3662 619112 3667 619168
rect -960 619110 3667 619112
rect -960 619020 480 619110
rect 3601 619107 3667 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580257 591018 580323 591021
rect 583520 591018 584960 591108
rect 580257 591016 584960 591018
rect 580257 590960 580262 591016
rect 580318 590960 584960 591016
rect 580257 590958 584960 590960
rect 580257 590955 580323 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3785 566946 3851 566949
rect -960 566944 3851 566946
rect -960 566888 3790 566944
rect 3846 566888 3851 566944
rect -960 566886 3851 566888
rect -960 566796 480 566886
rect 3785 566883 3851 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580349 537842 580415 537845
rect 583520 537842 584960 537932
rect 580349 537840 584960 537842
rect 580349 537784 580354 537840
rect 580410 537784 584960 537840
rect 580349 537782 584960 537784
rect 580349 537779 580415 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3325 527914 3391 527917
rect -960 527912 3391 527914
rect -960 527856 3330 527912
rect 3386 527856 3391 527912
rect -960 527854 3391 527856
rect -960 527764 480 527854
rect 3325 527851 3391 527854
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 579981 511322 580047 511325
rect 583520 511322 584960 511412
rect 579981 511320 584960 511322
rect 579981 511264 579986 511320
rect 580042 511264 584960 511320
rect 579981 511262 584960 511264
rect 579981 511259 580047 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3693 501802 3759 501805
rect -960 501800 3759 501802
rect -960 501744 3698 501800
rect 3754 501744 3759 501800
rect -960 501742 3759 501744
rect -960 501652 480 501742
rect 3693 501739 3759 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580441 484666 580507 484669
rect 583520 484666 584960 484756
rect 580441 484664 584960 484666
rect 580441 484608 580446 484664
rect 580502 484608 584960 484664
rect 580441 484606 584960 484608
rect 580441 484603 580507 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3877 475690 3943 475693
rect -960 475688 3943 475690
rect -960 475632 3882 475688
rect 3938 475632 3943 475688
rect -960 475630 3943 475632
rect -960 475540 480 475630
rect 3877 475627 3943 475630
rect 579613 471474 579679 471477
rect 583520 471474 584960 471564
rect 579613 471472 584960 471474
rect 579613 471416 579618 471472
rect 579674 471416 584960 471472
rect 579613 471414 584960 471416
rect 579613 471411 579679 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 579613 458146 579679 458149
rect 583520 458146 584960 458236
rect 579613 458144 584960 458146
rect 579613 458088 579618 458144
rect 579674 458088 584960 458144
rect 579613 458086 584960 458088
rect 579613 458083 579679 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 2957 449578 3023 449581
rect -960 449576 3023 449578
rect -960 449520 2962 449576
rect 3018 449520 3023 449576
rect -960 449518 3023 449520
rect -960 449428 480 449518
rect 2957 449515 3023 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580533 431626 580599 431629
rect 583520 431626 584960 431716
rect 580533 431624 584960 431626
rect 580533 431568 580538 431624
rect 580594 431568 584960 431624
rect 580533 431566 584960 431568
rect 580533 431563 580599 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580625 378450 580691 378453
rect 583520 378450 584960 378540
rect 580625 378448 584960 378450
rect 580625 378392 580630 378448
rect 580686 378392 584960 378448
rect 580625 378390 584960 378392
rect 580625 378387 580691 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3877 358458 3943 358461
rect -960 358456 3943 358458
rect -960 358400 3882 358456
rect 3938 358400 3943 358456
rect -960 358398 3943 358400
rect -960 358308 480 358398
rect 3877 358395 3943 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580717 325274 580783 325277
rect 583520 325274 584960 325364
rect 580717 325272 584960 325274
rect 580717 325216 580722 325272
rect 580778 325216 584960 325272
rect 580717 325214 584960 325216
rect 580717 325211 580783 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3141 319290 3207 319293
rect -960 319288 3207 319290
rect -960 319232 3146 319288
rect 3202 319232 3207 319288
rect -960 319230 3207 319232
rect -960 319140 480 319230
rect 3141 319227 3207 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3969 293178 4035 293181
rect -960 293176 4035 293178
rect -960 293120 3974 293176
rect 4030 293120 4035 293176
rect -960 293118 4035 293120
rect -960 293028 480 293118
rect 3969 293115 4035 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580809 272234 580875 272237
rect 583520 272234 584960 272324
rect 580809 272232 584960 272234
rect 580809 272176 580814 272232
rect 580870 272176 584960 272232
rect 580809 272174 584960 272176
rect 580809 272171 580875 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2865 254146 2931 254149
rect -960 254144 2931 254146
rect -960 254088 2870 254144
rect 2926 254088 2931 254144
rect -960 254086 2931 254088
rect -960 253996 480 254086
rect 2865 254083 2931 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 4061 241090 4127 241093
rect -960 241088 4127 241090
rect -960 241032 4066 241088
rect 4122 241032 4127 241088
rect -960 241030 4127 241032
rect -960 240940 480 241030
rect 4061 241027 4127 241030
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 579981 219058 580047 219061
rect 583520 219058 584960 219148
rect 579981 219056 584960 219058
rect 579981 219000 579986 219056
rect 580042 219000 584960 219056
rect 579981 218998 584960 219000
rect 579981 218995 580047 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 117313 137594 117379 137597
rect 117313 137592 120060 137594
rect 117313 137536 117318 137592
rect 117374 137536 120060 137592
rect 117313 137534 120060 137536
rect 117313 137531 117379 137534
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 117313 136098 117379 136101
rect 117313 136096 120060 136098
rect 117313 136040 117318 136096
rect 117374 136040 120060 136096
rect 117313 136038 120060 136040
rect 117313 136035 117379 136038
rect 117313 134602 117379 134605
rect 117313 134600 120060 134602
rect 117313 134544 117318 134600
rect 117374 134544 120060 134600
rect 117313 134542 120060 134544
rect 117313 134539 117379 134542
rect 117405 133106 117471 133109
rect 117405 133104 120060 133106
rect 117405 133048 117410 133104
rect 117466 133048 120060 133104
rect 117405 133046 120060 133048
rect 117405 133043 117471 133046
rect 117313 131610 117379 131613
rect 117313 131608 120060 131610
rect 117313 131552 117318 131608
rect 117374 131552 120060 131608
rect 117313 131550 120060 131552
rect 117313 131547 117379 131550
rect 189582 130525 189642 131036
rect 189582 130520 189691 130525
rect 189582 130464 189630 130520
rect 189686 130464 189691 130520
rect 189582 130462 189691 130464
rect 189625 130459 189691 130462
rect 117313 130114 117379 130117
rect 117313 130112 120060 130114
rect 117313 130056 117318 130112
rect 117374 130056 120060 130112
rect 117313 130054 120060 130056
rect 117313 130051 117379 130054
rect 190729 129706 190795 129709
rect 189796 129704 190795 129706
rect 189796 129648 190734 129704
rect 190790 129648 190795 129704
rect 189796 129646 190795 129648
rect 190729 129643 190795 129646
rect 117313 128618 117379 128621
rect 117313 128616 120060 128618
rect 117313 128560 117318 128616
rect 117374 128560 120060 128616
rect 117313 128558 120060 128560
rect 117313 128555 117379 128558
rect 191925 128346 191991 128349
rect 189796 128344 191991 128346
rect 189796 128288 191930 128344
rect 191986 128288 191991 128344
rect 189796 128286 191991 128288
rect 191925 128283 191991 128286
rect 117313 127122 117379 127125
rect 117313 127120 120060 127122
rect 117313 127064 117318 127120
rect 117374 127064 120060 127120
rect 117313 127062 120060 127064
rect 117313 127059 117379 127062
rect 191189 126986 191255 126989
rect 189796 126984 191255 126986
rect 189796 126928 191194 126984
rect 191250 126928 191255 126984
rect 189796 126926 191255 126928
rect 191189 126923 191255 126926
rect 189625 126170 189691 126173
rect 189582 126168 189691 126170
rect 189582 126112 189630 126168
rect 189686 126112 189691 126168
rect 189582 126107 189691 126112
rect 117313 125626 117379 125629
rect 117313 125624 120060 125626
rect 117313 125568 117318 125624
rect 117374 125568 120060 125624
rect 189582 125596 189642 126107
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 583520 125884 584960 125974
rect 117313 125566 120060 125568
rect 117313 125563 117379 125566
rect 190637 124266 190703 124269
rect 189796 124264 190703 124266
rect 189796 124208 190642 124264
rect 190698 124208 190703 124264
rect 189796 124206 190703 124208
rect 190637 124203 190703 124206
rect 117313 124130 117379 124133
rect 117313 124128 120060 124130
rect 117313 124072 117318 124128
rect 117374 124072 120060 124128
rect 117313 124070 120060 124072
rect 117313 124067 117379 124070
rect -960 123572 480 123812
rect 192017 122906 192083 122909
rect 189796 122904 192083 122906
rect 189796 122848 192022 122904
rect 192078 122848 192083 122904
rect 189796 122846 192083 122848
rect 192017 122843 192083 122846
rect 117313 122634 117379 122637
rect 117313 122632 120060 122634
rect 117313 122576 117318 122632
rect 117374 122576 120060 122632
rect 117313 122574 120060 122576
rect 117313 122571 117379 122574
rect 191097 121546 191163 121549
rect 189796 121544 191163 121546
rect 189796 121488 191102 121544
rect 191158 121488 191163 121544
rect 189796 121486 191163 121488
rect 191097 121483 191163 121486
rect 117313 121138 117379 121141
rect 117313 121136 120060 121138
rect 117313 121080 117318 121136
rect 117374 121080 120060 121136
rect 117313 121078 120060 121080
rect 117313 121075 117379 121078
rect 189349 120730 189415 120733
rect 189349 120728 189458 120730
rect 189349 120672 189354 120728
rect 189410 120672 189458 120728
rect 189349 120667 189458 120672
rect 189398 120156 189458 120667
rect 117313 119642 117379 119645
rect 117313 119640 120060 119642
rect 117313 119584 117318 119640
rect 117374 119584 120060 119640
rect 117313 119582 120060 119584
rect 117313 119579 117379 119582
rect 189717 119370 189783 119373
rect 189717 119368 189826 119370
rect 189717 119312 189722 119368
rect 189778 119312 189826 119368
rect 189717 119307 189826 119312
rect 189766 118796 189826 119307
rect 117313 118146 117379 118149
rect 117313 118144 120060 118146
rect 117313 118088 117318 118144
rect 117374 118088 120060 118144
rect 117313 118086 120060 118088
rect 117313 118083 117379 118086
rect 190545 117466 190611 117469
rect 189796 117464 190611 117466
rect 189796 117408 190550 117464
rect 190606 117408 190611 117464
rect 189796 117406 190611 117408
rect 190545 117403 190611 117406
rect 117313 116650 117379 116653
rect 189349 116650 189415 116653
rect 117313 116648 120060 116650
rect 117313 116592 117318 116648
rect 117374 116592 120060 116648
rect 117313 116590 120060 116592
rect 189349 116648 189458 116650
rect 189349 116592 189354 116648
rect 189410 116592 189458 116648
rect 117313 116587 117379 116590
rect 189349 116587 189458 116592
rect 189398 116076 189458 116587
rect 117313 115154 117379 115157
rect 117313 115152 120060 115154
rect 117313 115096 117318 115152
rect 117374 115096 120060 115152
rect 117313 115094 120060 115096
rect 117313 115091 117379 115094
rect 190821 114746 190887 114749
rect 189796 114744 190887 114746
rect 189796 114688 190826 114744
rect 190882 114688 190887 114744
rect 189796 114686 190887 114688
rect 190821 114683 190887 114686
rect 189441 113930 189507 113933
rect 189398 113928 189507 113930
rect 189398 113872 189446 113928
rect 189502 113872 189507 113928
rect 189398 113867 189507 113872
rect 118049 113658 118115 113661
rect 118049 113656 120060 113658
rect 118049 113600 118054 113656
rect 118110 113600 120060 113656
rect 118049 113598 120060 113600
rect 118049 113595 118115 113598
rect 189398 113356 189458 113867
rect 580073 112842 580139 112845
rect 583520 112842 584960 112932
rect 580073 112840 584960 112842
rect 580073 112784 580078 112840
rect 580134 112784 584960 112840
rect 580073 112782 584960 112784
rect 580073 112779 580139 112782
rect 583520 112692 584960 112782
rect 189533 112570 189599 112573
rect 189533 112568 189642 112570
rect 189533 112512 189538 112568
rect 189594 112512 189642 112568
rect 189533 112507 189642 112512
rect 119245 112162 119311 112165
rect 119245 112160 120060 112162
rect 119245 112104 119250 112160
rect 119306 112104 120060 112160
rect 119245 112102 120060 112104
rect 119245 112099 119311 112102
rect 189582 111996 189642 112507
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 118969 110666 119035 110669
rect 191005 110666 191071 110669
rect 118969 110664 120060 110666
rect 118969 110608 118974 110664
rect 119030 110608 120060 110664
rect 118969 110606 120060 110608
rect 189796 110664 191071 110666
rect 189796 110608 191010 110664
rect 191066 110608 191071 110664
rect 189796 110606 191071 110608
rect 118969 110603 119035 110606
rect 191005 110603 191071 110606
rect 190913 109306 190979 109309
rect 189796 109304 190979 109306
rect 189796 109248 190918 109304
rect 190974 109248 190979 109304
rect 189796 109246 190979 109248
rect 190913 109243 190979 109246
rect 119061 109170 119127 109173
rect 119061 109168 120060 109170
rect 119061 109112 119066 109168
rect 119122 109112 120060 109168
rect 119061 109110 120060 109112
rect 119061 109107 119127 109110
rect 191925 107946 191991 107949
rect 189796 107944 191991 107946
rect 189796 107888 191930 107944
rect 191986 107888 191991 107944
rect 189796 107886 191991 107888
rect 191925 107883 191991 107886
rect 119153 107674 119219 107677
rect 119153 107672 120060 107674
rect 119153 107616 119158 107672
rect 119214 107616 120060 107672
rect 119153 107614 120060 107616
rect 119153 107611 119219 107614
rect 191925 106586 191991 106589
rect 189796 106584 191991 106586
rect 189796 106528 191930 106584
rect 191986 106528 191991 106584
rect 189796 106526 191991 106528
rect 191925 106523 191991 106526
rect 118877 106178 118943 106181
rect 118877 106176 120060 106178
rect 118877 106120 118882 106176
rect 118938 106120 120060 106176
rect 118877 106118 120060 106120
rect 118877 106115 118943 106118
rect 191925 105226 191991 105229
rect 189796 105224 191991 105226
rect 189796 105168 191930 105224
rect 191986 105168 191991 105224
rect 189796 105166 191991 105168
rect 191925 105163 191991 105166
rect 118785 104682 118851 104685
rect 118785 104680 120060 104682
rect 118785 104624 118790 104680
rect 118846 104624 120060 104680
rect 118785 104622 120060 104624
rect 118785 104619 118851 104622
rect 193121 103866 193187 103869
rect 189796 103864 193187 103866
rect 189796 103808 193126 103864
rect 193182 103808 193187 103864
rect 189796 103806 193187 103808
rect 193121 103803 193187 103806
rect 118693 103186 118759 103189
rect 118693 103184 120060 103186
rect 118693 103128 118698 103184
rect 118754 103128 120060 103184
rect 118693 103126 120060 103128
rect 118693 103123 118759 103126
rect 193121 102506 193187 102509
rect 189796 102504 193187 102506
rect 189796 102448 193126 102504
rect 193182 102448 193187 102504
rect 189796 102446 193187 102448
rect 193121 102443 193187 102446
rect 120717 102098 120783 102101
rect 120582 102096 120783 102098
rect 120582 102040 120722 102096
rect 120778 102040 120783 102096
rect 120582 102038 120783 102040
rect 120582 101660 120642 102038
rect 120717 102035 120783 102038
rect 191925 101146 191991 101149
rect 189796 101144 191991 101146
rect 189796 101088 191930 101144
rect 191986 101088 191991 101144
rect 189796 101086 191991 101088
rect 191925 101083 191991 101086
rect 120809 100738 120875 100741
rect 120582 100736 120875 100738
rect 120582 100680 120814 100736
rect 120870 100680 120875 100736
rect 120582 100678 120875 100680
rect 120582 100164 120642 100678
rect 120809 100675 120875 100678
rect 192385 99786 192451 99789
rect 189796 99784 192451 99786
rect 189796 99728 192390 99784
rect 192446 99728 192451 99784
rect 189796 99726 192451 99728
rect 192385 99723 192451 99726
rect 579981 99514 580047 99517
rect 583520 99514 584960 99604
rect 579981 99512 584960 99514
rect 579981 99456 579986 99512
rect 580042 99456 584960 99512
rect 579981 99454 584960 99456
rect 579981 99451 580047 99454
rect 583520 99364 584960 99454
rect 120901 98698 120967 98701
rect 120612 98696 120967 98698
rect 120612 98640 120906 98696
rect 120962 98640 120967 98696
rect 120612 98638 120967 98640
rect 120901 98635 120967 98638
rect 192109 98426 192175 98429
rect 189796 98424 192175 98426
rect 189796 98368 192114 98424
rect 192170 98368 192175 98424
rect 189796 98366 192175 98368
rect 192109 98363 192175 98366
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 120993 97202 121059 97205
rect 120612 97200 121059 97202
rect 120612 97144 120998 97200
rect 121054 97144 121059 97200
rect 120612 97142 121059 97144
rect 120993 97139 121059 97142
rect 192201 97066 192267 97069
rect 189796 97064 192267 97066
rect 189796 97008 192206 97064
rect 192262 97008 192267 97064
rect 189796 97006 192267 97008
rect 192201 97003 192267 97006
rect 118601 95706 118667 95709
rect 191925 95706 191991 95709
rect 118601 95704 120060 95706
rect 118601 95648 118606 95704
rect 118662 95648 120060 95704
rect 118601 95646 120060 95648
rect 189796 95704 191991 95706
rect 189796 95648 191930 95704
rect 191986 95648 191991 95704
rect 189796 95646 191991 95648
rect 118601 95643 118667 95646
rect 191925 95643 191991 95646
rect 193121 94346 193187 94349
rect 189796 94344 193187 94346
rect 189796 94288 193126 94344
rect 193182 94288 193187 94344
rect 189796 94286 193187 94288
rect 193121 94283 193187 94286
rect 118509 94210 118575 94213
rect 118509 94208 120060 94210
rect 118509 94152 118514 94208
rect 118570 94152 120060 94208
rect 118509 94150 120060 94152
rect 118509 94147 118575 94150
rect 192569 92986 192635 92989
rect 189796 92984 192635 92986
rect 189796 92928 192574 92984
rect 192630 92928 192635 92984
rect 189796 92926 192635 92928
rect 192569 92923 192635 92926
rect 118233 92714 118299 92717
rect 118233 92712 120060 92714
rect 118233 92656 118238 92712
rect 118294 92656 120060 92712
rect 118233 92654 120060 92656
rect 118233 92651 118299 92654
rect 193121 91626 193187 91629
rect 189796 91624 193187 91626
rect 189796 91568 193126 91624
rect 193182 91568 193187 91624
rect 189796 91566 193187 91568
rect 193121 91563 193187 91566
rect 118141 91218 118207 91221
rect 118141 91216 120060 91218
rect 118141 91160 118146 91216
rect 118202 91160 120060 91216
rect 118141 91158 120060 91160
rect 118141 91155 118207 91158
rect 193121 90266 193187 90269
rect 189796 90264 193187 90266
rect 189796 90208 193126 90264
rect 193182 90208 193187 90264
rect 189796 90206 193187 90208
rect 193121 90203 193187 90206
rect 118417 89722 118483 89725
rect 118417 89720 120060 89722
rect 118417 89664 118422 89720
rect 118478 89664 120060 89720
rect 118417 89662 120060 89664
rect 118417 89659 118483 89662
rect 193121 88906 193187 88909
rect 189796 88904 193187 88906
rect 189796 88848 193126 88904
rect 193182 88848 193187 88904
rect 189796 88846 193187 88848
rect 193121 88843 193187 88846
rect 118325 88226 118391 88229
rect 118325 88224 120060 88226
rect 118325 88168 118330 88224
rect 118386 88168 120060 88224
rect 118325 88166 120060 88168
rect 118325 88163 118391 88166
rect 192937 87546 193003 87549
rect 189796 87544 193003 87546
rect 189796 87488 192942 87544
rect 192998 87488 193003 87544
rect 189796 87486 193003 87488
rect 192937 87483 193003 87486
rect 118509 86730 118575 86733
rect 118509 86728 120060 86730
rect 118509 86672 118514 86728
rect 118570 86672 120060 86728
rect 118509 86670 120060 86672
rect 118509 86667 118575 86670
rect 193029 86186 193095 86189
rect 189796 86184 193095 86186
rect 189796 86128 193034 86184
rect 193090 86128 193095 86184
rect 189796 86126 193095 86128
rect 193029 86123 193095 86126
rect 580809 86186 580875 86189
rect 583520 86186 584960 86276
rect 580809 86184 584960 86186
rect 580809 86128 580814 86184
rect 580870 86128 584960 86184
rect 580809 86126 584960 86128
rect 580809 86123 580875 86126
rect 583520 86036 584960 86126
rect 118601 85234 118667 85237
rect 118601 85232 120060 85234
rect 118601 85176 118606 85232
rect 118662 85176 120060 85232
rect 118601 85174 120060 85176
rect 118601 85171 118667 85174
rect 193121 84826 193187 84829
rect 189796 84824 193187 84826
rect -960 84690 480 84780
rect 189796 84768 193126 84824
rect 193182 84768 193187 84824
rect 189796 84766 193187 84768
rect 193121 84763 193187 84766
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 118417 83738 118483 83741
rect 118417 83736 120060 83738
rect 118417 83680 118422 83736
rect 118478 83680 120060 83736
rect 118417 83678 120060 83680
rect 118417 83675 118483 83678
rect 193121 83466 193187 83469
rect 189796 83464 193187 83466
rect 189796 83408 193126 83464
rect 193182 83408 193187 83464
rect 189796 83406 193187 83408
rect 193121 83403 193187 83406
rect 189349 82378 189415 82381
rect 580390 82378 580396 82380
rect 189349 82376 580396 82378
rect 189349 82320 189354 82376
rect 189410 82320 580396 82376
rect 189349 82318 580396 82320
rect 189349 82315 189415 82318
rect 580390 82316 580396 82318
rect 580460 82316 580466 82380
rect 120582 81698 120642 82212
rect 192569 82106 192635 82109
rect 189796 82104 192635 82106
rect 189796 82048 192574 82104
rect 192630 82048 192635 82104
rect 189796 82046 192635 82048
rect 192569 82043 192635 82046
rect 120717 81698 120783 81701
rect 120582 81696 120783 81698
rect 120582 81640 120722 81696
rect 120778 81640 120783 81696
rect 120582 81638 120783 81640
rect 120717 81635 120783 81638
rect 193121 80746 193187 80749
rect 189796 80744 193187 80746
rect 189796 80688 193126 80744
rect 193182 80688 193187 80744
rect 189796 80686 193187 80688
rect 193121 80683 193187 80686
rect 118601 80610 118667 80613
rect 580809 80610 580875 80613
rect 118601 80608 580875 80610
rect 118601 80552 118606 80608
rect 118662 80552 580814 80608
rect 580870 80552 580875 80608
rect 118601 80550 580875 80552
rect 118601 80547 118667 80550
rect 580809 80547 580875 80550
rect 164366 80412 164372 80476
rect 164436 80474 164442 80476
rect 433333 80474 433399 80477
rect 164436 80472 433399 80474
rect 164436 80416 433338 80472
rect 433394 80416 433399 80472
rect 164436 80414 433399 80416
rect 164436 80412 164442 80414
rect 433333 80411 433399 80414
rect 177982 80338 177988 80340
rect 164190 80278 177988 80338
rect 140814 80140 140820 80204
rect 140884 80202 140890 80204
rect 140884 80142 143688 80202
rect 140884 80140 140890 80142
rect 134190 80004 134196 80068
rect 134260 80066 134266 80068
rect 134260 80006 134626 80066
rect 134260 80004 134266 80006
rect 131067 79962 131133 79967
rect 130101 79930 130167 79933
rect 131067 79930 131072 79962
rect 130101 79928 131072 79930
rect 130101 79872 130106 79928
rect 130162 79906 131072 79928
rect 131128 79906 131133 79962
rect 131435 79962 131501 79967
rect 130162 79901 131133 79906
rect 130162 79872 131130 79901
rect 130101 79870 131130 79872
rect 130101 79867 130167 79870
rect 131246 79868 131252 79932
rect 131316 79930 131322 79932
rect 131435 79930 131440 79962
rect 131316 79906 131440 79930
rect 131496 79906 131501 79962
rect 131316 79901 131501 79906
rect 131803 79962 131869 79967
rect 131803 79906 131808 79962
rect 131864 79906 131869 79962
rect 132171 79962 132237 79967
rect 131803 79901 131869 79906
rect 131316 79870 131498 79901
rect 131316 79868 131322 79870
rect 131806 79797 131866 79901
rect 131982 79868 131988 79932
rect 132052 79930 132058 79932
rect 132171 79930 132176 79962
rect 132052 79906 132176 79930
rect 132232 79906 132237 79962
rect 132355 79962 132421 79967
rect 132355 79932 132360 79962
rect 132416 79932 132421 79962
rect 132907 79962 132973 79967
rect 132052 79901 132237 79906
rect 132052 79870 132234 79901
rect 132052 79868 132058 79870
rect 132350 79868 132356 79932
rect 132420 79930 132426 79932
rect 132723 79930 132789 79933
rect 132907 79932 132912 79962
rect 132968 79932 132973 79962
rect 133275 79962 133341 79967
rect 132420 79870 132478 79930
rect 132542 79928 132789 79930
rect 132542 79872 132728 79928
rect 132784 79872 132789 79928
rect 132542 79870 132789 79872
rect 132420 79868 132426 79870
rect 131757 79792 131866 79797
rect 131757 79736 131762 79792
rect 131818 79736 131866 79792
rect 131757 79734 131866 79736
rect 132217 79794 132283 79797
rect 132542 79794 132602 79870
rect 132723 79867 132789 79870
rect 132902 79868 132908 79932
rect 132972 79930 132978 79932
rect 132972 79870 133030 79930
rect 133275 79906 133280 79962
rect 133336 79906 133341 79962
rect 133643 79962 133709 79967
rect 133275 79901 133341 79906
rect 133459 79928 133525 79933
rect 132972 79868 132978 79870
rect 133278 79797 133338 79901
rect 133459 79872 133464 79928
rect 133520 79872 133525 79928
rect 133643 79906 133648 79962
rect 133704 79906 133709 79962
rect 133643 79901 133709 79906
rect 134011 79962 134077 79967
rect 134011 79906 134016 79962
rect 134072 79930 134077 79962
rect 134374 79930 134380 79932
rect 134072 79906 134380 79930
rect 134011 79901 134380 79906
rect 133459 79867 133525 79872
rect 133462 79797 133522 79867
rect 133646 79797 133706 79901
rect 134014 79870 134380 79901
rect 134374 79868 134380 79870
rect 134444 79868 134450 79932
rect 132217 79792 132602 79794
rect 132217 79736 132222 79792
rect 132278 79736 132602 79792
rect 132217 79734 132602 79736
rect 132677 79794 132743 79797
rect 133086 79794 133092 79796
rect 132677 79792 133092 79794
rect 132677 79736 132682 79792
rect 132738 79736 133092 79792
rect 132677 79734 133092 79736
rect 131757 79731 131823 79734
rect 132217 79731 132283 79734
rect 132677 79731 132743 79734
rect 133086 79732 133092 79734
rect 133156 79732 133162 79796
rect 133229 79792 133338 79797
rect 133229 79736 133234 79792
rect 133290 79736 133338 79792
rect 133229 79734 133338 79736
rect 133413 79792 133522 79797
rect 133413 79736 133418 79792
rect 133474 79736 133522 79792
rect 133413 79734 133522 79736
rect 133597 79792 133706 79797
rect 133597 79736 133602 79792
rect 133658 79736 133706 79792
rect 133597 79734 133706 79736
rect 134057 79794 134123 79797
rect 134190 79794 134196 79796
rect 134057 79792 134196 79794
rect 134057 79736 134062 79792
rect 134118 79736 134196 79792
rect 134057 79734 134196 79736
rect 133229 79731 133295 79734
rect 133413 79731 133479 79734
rect 133597 79731 133663 79734
rect 134057 79731 134123 79734
rect 134190 79732 134196 79734
rect 134260 79732 134266 79796
rect 134379 79794 134445 79797
rect 134566 79794 134626 80006
rect 143206 80004 143212 80068
rect 143276 80066 143282 80068
rect 143276 80006 143550 80066
rect 143276 80004 143282 80006
rect 138335 79964 138401 79967
rect 139623 79964 139689 79967
rect 138335 79962 138444 79964
rect 135023 79930 135089 79933
rect 134379 79792 134626 79794
rect 134379 79736 134384 79792
rect 134440 79736 134626 79792
rect 134379 79734 134626 79736
rect 134796 79928 135089 79930
rect 134796 79872 135028 79928
rect 135084 79872 135089 79928
rect 134796 79870 135089 79872
rect 134796 79794 134856 79870
rect 135023 79867 135089 79870
rect 135294 79868 135300 79932
rect 135364 79930 135370 79932
rect 135483 79930 135549 79933
rect 135364 79928 135549 79930
rect 135364 79872 135488 79928
rect 135544 79872 135549 79928
rect 135364 79870 135549 79872
rect 135364 79868 135370 79870
rect 135483 79867 135549 79870
rect 136214 79868 136220 79932
rect 136284 79930 136290 79932
rect 136495 79930 136561 79933
rect 136284 79928 136561 79930
rect 136284 79872 136500 79928
rect 136556 79872 136561 79928
rect 136284 79870 136561 79872
rect 136284 79868 136290 79870
rect 136495 79867 136561 79870
rect 137047 79930 137113 79933
rect 137686 79930 137692 79932
rect 137047 79928 137692 79930
rect 137047 79872 137052 79928
rect 137108 79872 137692 79928
rect 137047 79870 137692 79872
rect 137047 79867 137113 79870
rect 137686 79868 137692 79870
rect 137756 79868 137762 79932
rect 137870 79868 137876 79932
rect 137940 79930 137946 79932
rect 138335 79930 138340 79962
rect 137940 79906 138340 79930
rect 138396 79906 138444 79962
rect 139488 79962 139689 79964
rect 137940 79870 138444 79906
rect 138519 79930 138585 79933
rect 138979 79932 139045 79933
rect 138519 79928 138858 79930
rect 138519 79872 138524 79928
rect 138580 79872 138858 79928
rect 138519 79870 138858 79872
rect 137940 79868 137946 79870
rect 138519 79867 138585 79870
rect 134926 79794 134932 79796
rect 134796 79734 134932 79794
rect 134379 79731 134445 79734
rect 134926 79732 134932 79734
rect 134996 79732 135002 79796
rect 135253 79794 135319 79797
rect 135478 79794 135484 79796
rect 135253 79792 135484 79794
rect 135253 79736 135258 79792
rect 135314 79736 135484 79792
rect 135253 79734 135484 79736
rect 135253 79731 135319 79734
rect 135478 79732 135484 79734
rect 135548 79732 135554 79796
rect 135667 79794 135733 79797
rect 135846 79794 135852 79796
rect 135667 79792 135852 79794
rect 135667 79736 135672 79792
rect 135728 79736 135852 79792
rect 135667 79734 135852 79736
rect 135667 79731 135733 79734
rect 135846 79732 135852 79734
rect 135916 79732 135922 79796
rect 136633 79794 136699 79797
rect 137139 79794 137205 79797
rect 136633 79792 137205 79794
rect 136633 79736 136638 79792
rect 136694 79736 137144 79792
rect 137200 79736 137205 79792
rect 136633 79734 137205 79736
rect 136633 79731 136699 79734
rect 137139 79731 137205 79734
rect 138289 79794 138355 79797
rect 138422 79794 138428 79796
rect 138289 79792 138428 79794
rect 138289 79736 138294 79792
rect 138350 79736 138428 79792
rect 138289 79734 138428 79736
rect 138289 79731 138355 79734
rect 138422 79732 138428 79734
rect 138492 79732 138498 79796
rect 138798 79794 138858 79870
rect 138974 79868 138980 79932
rect 139044 79930 139050 79932
rect 139044 79870 139136 79930
rect 139044 79868 139050 79870
rect 139342 79868 139348 79932
rect 139412 79930 139418 79932
rect 139488 79930 139628 79962
rect 139412 79906 139628 79930
rect 139684 79906 139689 79962
rect 140267 79962 140333 79967
rect 139412 79904 139689 79906
rect 139412 79870 139548 79904
rect 139623 79901 139689 79904
rect 139899 79928 139965 79933
rect 139899 79872 139904 79928
rect 139960 79872 139965 79928
rect 140267 79906 140272 79962
rect 140328 79906 140333 79962
rect 143490 79933 143550 80006
rect 143628 79967 143688 80142
rect 148358 80140 148364 80204
rect 148428 80202 148434 80204
rect 148428 80142 148886 80202
rect 148428 80140 148434 80142
rect 143628 79962 143737 79967
rect 140267 79901 140333 79906
rect 140727 79928 140793 79933
rect 139412 79868 139418 79870
rect 138979 79867 139045 79868
rect 139899 79867 139965 79872
rect 138933 79794 138999 79797
rect 138798 79792 138999 79794
rect 138798 79736 138938 79792
rect 138994 79736 138999 79792
rect 138798 79734 138999 79736
rect 138933 79731 138999 79734
rect 139710 79732 139716 79796
rect 139780 79794 139786 79796
rect 139902 79794 139962 79867
rect 139780 79734 139962 79794
rect 140129 79794 140195 79797
rect 140270 79794 140330 79901
rect 140727 79872 140732 79928
rect 140788 79872 140793 79928
rect 140727 79867 140793 79872
rect 141366 79868 141372 79932
rect 141436 79930 141442 79932
rect 141647 79930 141713 79933
rect 142659 79932 142725 79933
rect 142654 79930 142660 79932
rect 141436 79928 141713 79930
rect 141436 79872 141652 79928
rect 141708 79872 141713 79928
rect 141436 79870 141713 79872
rect 142568 79870 142660 79930
rect 141436 79868 141442 79870
rect 141647 79867 141713 79870
rect 142654 79868 142660 79870
rect 142724 79868 142730 79932
rect 143487 79928 143553 79933
rect 143487 79872 143492 79928
rect 143548 79872 143553 79928
rect 143628 79906 143676 79962
rect 143732 79906 143737 79962
rect 147443 79962 147509 79967
rect 143628 79904 143737 79906
rect 143671 79901 143737 79904
rect 142659 79867 142725 79868
rect 143487 79867 143553 79872
rect 143942 79868 143948 79932
rect 144012 79930 144018 79932
rect 144223 79930 144289 79933
rect 144683 79932 144749 79933
rect 144678 79930 144684 79932
rect 144012 79928 144289 79930
rect 144012 79872 144228 79928
rect 144284 79872 144289 79928
rect 144012 79870 144289 79872
rect 144592 79870 144684 79930
rect 144012 79868 144018 79870
rect 144223 79867 144289 79870
rect 144678 79868 144684 79870
rect 144748 79868 144754 79932
rect 145230 79868 145236 79932
rect 145300 79930 145306 79932
rect 145879 79930 145945 79933
rect 145300 79928 145945 79930
rect 145300 79872 145884 79928
rect 145940 79872 145945 79928
rect 145300 79870 145945 79872
rect 145300 79868 145306 79870
rect 144683 79867 144749 79868
rect 145879 79867 145945 79870
rect 146886 79868 146892 79932
rect 146956 79930 146962 79932
rect 147075 79930 147141 79933
rect 146956 79928 147141 79930
rect 146956 79872 147080 79928
rect 147136 79872 147141 79928
rect 147443 79906 147448 79962
rect 147504 79906 147509 79962
rect 148455 79962 148521 79967
rect 147443 79901 147509 79906
rect 146956 79870 147141 79872
rect 146956 79868 146962 79870
rect 147075 79867 147141 79870
rect 140129 79792 140330 79794
rect 140129 79736 140134 79792
rect 140190 79736 140330 79792
rect 140129 79734 140330 79736
rect 140589 79794 140655 79797
rect 140730 79794 140790 79867
rect 141187 79826 141253 79831
rect 140589 79792 140790 79794
rect 140589 79736 140594 79792
rect 140650 79736 140790 79792
rect 140589 79734 140790 79736
rect 139780 79732 139786 79734
rect 140129 79731 140195 79734
rect 140589 79731 140655 79734
rect 140998 79732 141004 79796
rect 141068 79794 141074 79796
rect 141187 79794 141192 79826
rect 141068 79770 141192 79794
rect 141248 79770 141253 79826
rect 143441 79796 143507 79797
rect 143390 79794 143396 79796
rect 141068 79765 141253 79770
rect 141068 79734 141250 79765
rect 143350 79734 143396 79794
rect 143460 79792 143507 79796
rect 143502 79736 143507 79792
rect 141068 79732 141074 79734
rect 143390 79732 143396 79734
rect 143460 79732 143507 79736
rect 144126 79732 144132 79796
rect 144196 79794 144202 79796
rect 144821 79794 144887 79797
rect 146523 79796 146589 79797
rect 146518 79794 146524 79796
rect 144196 79792 144887 79794
rect 144196 79736 144826 79792
rect 144882 79736 144887 79792
rect 144196 79734 144887 79736
rect 146432 79734 146524 79794
rect 144196 79732 144202 79734
rect 143441 79731 143507 79732
rect 144821 79731 144887 79734
rect 146518 79732 146524 79734
rect 146588 79732 146594 79796
rect 147070 79732 147076 79796
rect 147140 79794 147146 79796
rect 147446 79794 147506 79901
rect 148174 79868 148180 79932
rect 148244 79930 148250 79932
rect 148455 79930 148460 79962
rect 148244 79906 148460 79930
rect 148516 79906 148521 79962
rect 148244 79901 148521 79906
rect 148639 79964 148705 79967
rect 148639 79962 148748 79964
rect 148639 79906 148644 79962
rect 148700 79906 148748 79962
rect 148826 79933 148886 80142
rect 151302 80140 151308 80204
rect 151372 80202 151378 80204
rect 164190 80202 164250 80278
rect 177982 80276 177988 80278
rect 178052 80276 178058 80340
rect 151372 80142 153486 80202
rect 151372 80140 151378 80142
rect 153426 79967 153486 80142
rect 157382 80142 164250 80202
rect 149099 79962 149165 79967
rect 149559 79964 149625 79967
rect 148639 79901 148748 79906
rect 148244 79870 148518 79901
rect 148244 79868 148250 79870
rect 147140 79734 147506 79794
rect 148688 79796 148748 79901
rect 148823 79928 148889 79933
rect 149099 79932 149104 79962
rect 149160 79932 149165 79962
rect 149516 79962 149625 79964
rect 149516 79932 149564 79962
rect 148823 79872 148828 79928
rect 148884 79872 148889 79928
rect 148823 79867 148889 79872
rect 149094 79868 149100 79932
rect 149164 79930 149170 79932
rect 149164 79870 149222 79930
rect 149164 79868 149170 79870
rect 149462 79868 149468 79932
rect 149532 79906 149564 79932
rect 149620 79906 149625 79962
rect 150295 79962 150361 79967
rect 149743 79930 149809 79933
rect 149532 79901 149625 79906
rect 149700 79928 149809 79930
rect 149532 79870 149576 79901
rect 149700 79872 149748 79928
rect 149804 79872 149809 79928
rect 150295 79906 150300 79962
rect 150356 79906 150361 79962
rect 150755 79962 150821 79967
rect 150755 79932 150760 79962
rect 150816 79932 150821 79962
rect 150939 79962 151005 79967
rect 150295 79901 150361 79906
rect 149532 79868 149538 79870
rect 149700 79867 149809 79872
rect 148688 79734 148732 79796
rect 147140 79732 147146 79734
rect 148726 79732 148732 79734
rect 148796 79732 148802 79796
rect 149053 79794 149119 79797
rect 149700 79794 149760 79867
rect 149053 79792 149760 79794
rect 149053 79736 149058 79792
rect 149114 79736 149760 79792
rect 149053 79734 149760 79736
rect 146523 79731 146589 79732
rect 149053 79731 149119 79734
rect 149830 79732 149836 79796
rect 149900 79794 149906 79796
rect 150298 79794 150358 79901
rect 150750 79868 150756 79932
rect 150820 79930 150826 79932
rect 150820 79870 150878 79930
rect 150939 79906 150944 79962
rect 151000 79930 151005 79962
rect 151675 79962 151741 79967
rect 152319 79964 152385 79967
rect 151675 79932 151680 79962
rect 151736 79932 151741 79962
rect 152276 79962 152385 79964
rect 152276 79932 152324 79962
rect 151118 79930 151124 79932
rect 151000 79906 151124 79930
rect 150939 79901 151124 79906
rect 150942 79870 151124 79901
rect 150820 79868 150826 79870
rect 151118 79868 151124 79870
rect 151188 79868 151194 79932
rect 151670 79868 151676 79932
rect 151740 79930 151746 79932
rect 151740 79870 151798 79930
rect 151740 79868 151746 79870
rect 152222 79868 152228 79932
rect 152292 79906 152324 79932
rect 152380 79906 152385 79962
rect 152871 79964 152937 79967
rect 152871 79962 152980 79964
rect 152292 79901 152385 79906
rect 152687 79930 152753 79933
rect 152687 79928 152796 79930
rect 152292 79870 152336 79901
rect 152687 79872 152692 79928
rect 152748 79872 152796 79928
rect 152871 79906 152876 79962
rect 152932 79932 152980 79962
rect 153423 79962 153489 79967
rect 152932 79906 152964 79932
rect 152871 79901 152964 79906
rect 152292 79868 152298 79870
rect 152687 79867 152796 79872
rect 152920 79870 152964 79901
rect 152958 79868 152964 79870
rect 153028 79868 153034 79932
rect 153423 79906 153428 79962
rect 153484 79906 153489 79962
rect 154435 79962 154501 79967
rect 153699 79932 153765 79933
rect 153694 79930 153700 79932
rect 153423 79901 153489 79906
rect 153608 79870 153700 79930
rect 153694 79868 153700 79870
rect 153764 79868 153770 79932
rect 154062 79868 154068 79932
rect 154132 79930 154138 79932
rect 154435 79930 154440 79962
rect 154132 79906 154440 79930
rect 154496 79906 154501 79962
rect 155355 79962 155421 79967
rect 154132 79901 154501 79906
rect 154132 79870 154498 79901
rect 154132 79868 154138 79870
rect 154614 79868 154620 79932
rect 154684 79930 154690 79932
rect 154895 79930 154961 79933
rect 154684 79928 154961 79930
rect 154684 79872 154900 79928
rect 154956 79872 154961 79928
rect 155355 79906 155360 79962
rect 155416 79906 155421 79962
rect 155539 79962 155605 79967
rect 155539 79932 155544 79962
rect 155600 79932 155605 79962
rect 155815 79964 155881 79967
rect 155815 79962 155924 79964
rect 155355 79901 155421 79906
rect 154684 79870 154961 79872
rect 154684 79868 154690 79870
rect 153699 79867 153765 79868
rect 154895 79867 154961 79870
rect 149900 79734 150358 79794
rect 149900 79732 149906 79734
rect 152406 79732 152412 79796
rect 152476 79794 152482 79796
rect 152736 79794 152796 79867
rect 155358 79797 155418 79901
rect 155534 79868 155540 79932
rect 155604 79930 155610 79932
rect 155604 79870 155662 79930
rect 155815 79906 155820 79962
rect 155876 79932 155924 79962
rect 156459 79962 156525 79967
rect 156459 79932 156464 79962
rect 156520 79932 156525 79962
rect 155876 79906 155908 79932
rect 155815 79901 155908 79906
rect 155864 79870 155908 79901
rect 155604 79868 155610 79870
rect 155902 79868 155908 79870
rect 155972 79868 155978 79932
rect 156454 79868 156460 79932
rect 156524 79930 156530 79932
rect 156735 79930 156801 79933
rect 157006 79930 157012 79932
rect 156524 79870 156582 79930
rect 156735 79928 157012 79930
rect 156735 79872 156740 79928
rect 156796 79872 157012 79928
rect 156735 79870 157012 79872
rect 156524 79868 156530 79870
rect 156735 79867 156801 79870
rect 157006 79868 157012 79870
rect 157076 79868 157082 79932
rect 152476 79734 152796 79794
rect 155309 79792 155418 79797
rect 156643 79796 156709 79797
rect 156638 79794 156644 79796
rect 155309 79736 155314 79792
rect 155370 79736 155418 79792
rect 155309 79734 155418 79736
rect 156552 79734 156644 79794
rect 152476 79732 152482 79734
rect 155309 79731 155375 79734
rect 156638 79732 156644 79734
rect 156708 79732 156714 79796
rect 156822 79732 156828 79796
rect 156892 79794 156898 79796
rect 157011 79794 157077 79797
rect 156892 79792 157077 79794
rect 156892 79736 157016 79792
rect 157072 79736 157077 79792
rect 156892 79734 157077 79736
rect 156892 79732 156898 79734
rect 156643 79731 156709 79732
rect 157011 79731 157077 79734
rect 6913 79658 6979 79661
rect 157382 79658 157442 80142
rect 168598 80140 168604 80204
rect 168668 80202 168674 80204
rect 168668 80142 179154 80202
rect 168668 80140 168674 80142
rect 163814 80004 163820 80068
rect 163884 80004 163890 80068
rect 171358 80004 171364 80068
rect 171428 80066 171434 80068
rect 171428 80004 171472 80066
rect 174302 80004 174308 80068
rect 174372 80066 174378 80068
rect 177062 80066 177068 80068
rect 174372 80006 174876 80066
rect 174372 80004 174378 80006
rect 157747 79962 157813 79967
rect 157747 79906 157752 79962
rect 157808 79906 157813 79962
rect 157931 79962 157997 79967
rect 157931 79932 157936 79962
rect 157992 79932 157997 79962
rect 160507 79962 160573 79967
rect 161335 79964 161401 79967
rect 157747 79901 157813 79906
rect 157750 79661 157810 79901
rect 157926 79868 157932 79932
rect 157996 79930 158002 79932
rect 157996 79870 158054 79930
rect 157996 79868 158002 79870
rect 158294 79868 158300 79932
rect 158364 79930 158370 79932
rect 158483 79930 158549 79933
rect 158364 79928 158549 79930
rect 158364 79872 158488 79928
rect 158544 79872 158549 79928
rect 158364 79870 158549 79872
rect 158364 79868 158370 79870
rect 158483 79867 158549 79870
rect 159311 79930 159377 79933
rect 160507 79932 160512 79962
rect 160568 79932 160573 79962
rect 161292 79962 161401 79964
rect 159311 79928 160202 79930
rect 159311 79872 159316 79928
rect 159372 79872 160202 79928
rect 159311 79870 160202 79872
rect 159311 79867 159377 79870
rect 158110 79732 158116 79796
rect 158180 79794 158186 79796
rect 158575 79794 158641 79797
rect 158180 79792 158641 79794
rect 158180 79736 158580 79792
rect 158636 79736 158641 79792
rect 158180 79734 158641 79736
rect 158180 79732 158186 79734
rect 158575 79731 158641 79734
rect 6913 79656 157442 79658
rect 6913 79600 6918 79656
rect 6974 79600 157442 79656
rect 6913 79598 157442 79600
rect 157701 79656 157810 79661
rect 157701 79600 157706 79656
rect 157762 79600 157810 79656
rect 157701 79598 157810 79600
rect 158345 79658 158411 79661
rect 158478 79658 158484 79660
rect 158345 79656 158484 79658
rect 158345 79600 158350 79656
rect 158406 79600 158484 79656
rect 158345 79598 158484 79600
rect 6913 79595 6979 79598
rect 157701 79595 157767 79598
rect 158345 79595 158411 79598
rect 158478 79596 158484 79598
rect 158548 79596 158554 79660
rect 159265 79658 159331 79661
rect 159633 79658 159699 79661
rect 159265 79656 159699 79658
rect 159265 79600 159270 79656
rect 159326 79600 159638 79656
rect 159694 79600 159699 79656
rect 159265 79598 159699 79600
rect 160142 79658 160202 79870
rect 160502 79868 160508 79932
rect 160572 79930 160578 79932
rect 160967 79930 161033 79933
rect 161292 79932 161340 79962
rect 160572 79870 160630 79930
rect 160967 79928 161168 79930
rect 160967 79872 160972 79928
rect 161028 79872 161168 79928
rect 160967 79870 161168 79872
rect 160572 79868 160578 79870
rect 160967 79867 161033 79870
rect 161108 79797 161168 79870
rect 161238 79868 161244 79932
rect 161308 79906 161340 79932
rect 161396 79906 161401 79962
rect 161979 79962 162045 79967
rect 161611 79932 161677 79933
rect 161979 79932 161984 79962
rect 162040 79932 162045 79962
rect 162347 79962 162413 79967
rect 162347 79932 162352 79962
rect 162408 79932 162413 79962
rect 162715 79962 162781 79967
rect 162715 79932 162720 79962
rect 162776 79932 162781 79962
rect 163635 79962 163701 79967
rect 161606 79930 161612 79932
rect 161308 79901 161401 79906
rect 161308 79870 161352 79901
rect 161520 79870 161612 79930
rect 161308 79868 161314 79870
rect 161606 79868 161612 79870
rect 161676 79868 161682 79932
rect 161974 79868 161980 79932
rect 162044 79930 162050 79932
rect 162044 79870 162102 79930
rect 162044 79868 162050 79870
rect 162342 79868 162348 79932
rect 162412 79930 162418 79932
rect 162412 79870 162470 79930
rect 162412 79868 162418 79870
rect 162710 79868 162716 79932
rect 162780 79930 162786 79932
rect 163175 79930 163241 79933
rect 163635 79932 163640 79962
rect 163696 79932 163701 79962
rect 162780 79870 162838 79930
rect 163175 79928 163514 79930
rect 163175 79872 163180 79928
rect 163236 79872 163514 79928
rect 163175 79870 163514 79872
rect 162780 79868 162786 79870
rect 161611 79867 161677 79868
rect 163175 79867 163241 79870
rect 161105 79792 161171 79797
rect 161105 79736 161110 79792
rect 161166 79736 161171 79792
rect 161105 79731 161171 79736
rect 162439 79794 162505 79797
rect 163454 79794 163514 79870
rect 163630 79868 163636 79932
rect 163700 79930 163706 79932
rect 163822 79930 163882 80004
rect 164371 79962 164437 79967
rect 164095 79930 164161 79933
rect 164371 79932 164376 79962
rect 164432 79932 164437 79962
rect 167683 79962 167749 79967
rect 163700 79870 163758 79930
rect 163822 79928 164161 79930
rect 163822 79872 164100 79928
rect 164156 79872 164161 79928
rect 163822 79870 164161 79872
rect 163700 79868 163706 79870
rect 164095 79867 164161 79870
rect 164366 79868 164372 79932
rect 164436 79930 164442 79932
rect 164739 79930 164805 79933
rect 164436 79870 164494 79930
rect 164558 79928 164805 79930
rect 164558 79872 164744 79928
rect 164800 79872 164805 79928
rect 164558 79870 164805 79872
rect 164436 79868 164442 79870
rect 163998 79794 164004 79796
rect 162439 79792 162548 79794
rect 162439 79736 162444 79792
rect 162500 79736 162548 79792
rect 162439 79731 162548 79736
rect 163454 79734 164004 79794
rect 163998 79732 164004 79734
rect 164068 79732 164074 79796
rect 161197 79658 161263 79661
rect 160142 79656 161263 79658
rect 160142 79600 161202 79656
rect 161258 79600 161263 79656
rect 160142 79598 161263 79600
rect 162488 79660 162548 79731
rect 164558 79661 164618 79870
rect 164739 79867 164805 79870
rect 164918 79868 164924 79932
rect 164988 79930 164994 79932
rect 165199 79930 165265 79933
rect 164988 79928 165265 79930
rect 164988 79872 165204 79928
rect 165260 79872 165265 79928
rect 164988 79870 165265 79872
rect 164988 79868 164994 79870
rect 165199 79867 165265 79870
rect 165475 79928 165541 79933
rect 166579 79932 166645 79933
rect 166574 79930 166580 79932
rect 165475 79872 165480 79928
rect 165536 79872 165541 79928
rect 165475 79867 165541 79872
rect 166488 79870 166580 79930
rect 166574 79868 166580 79870
rect 166644 79868 166650 79932
rect 166758 79868 166764 79932
rect 166828 79930 166834 79932
rect 167039 79930 167105 79933
rect 166828 79928 167105 79930
rect 166828 79872 167044 79928
rect 167100 79872 167105 79928
rect 166828 79870 167105 79872
rect 166828 79868 166834 79870
rect 166579 79867 166645 79868
rect 167039 79867 167105 79870
rect 167310 79868 167316 79932
rect 167380 79930 167386 79932
rect 167499 79930 167565 79933
rect 167380 79928 167565 79930
rect 167380 79872 167504 79928
rect 167560 79872 167565 79928
rect 167683 79906 167688 79962
rect 167744 79906 167749 79962
rect 168327 79962 168393 79967
rect 167683 79901 167749 79906
rect 167380 79870 167565 79872
rect 167380 79868 167386 79870
rect 167499 79867 167565 79870
rect 162488 79598 162532 79660
rect 159265 79595 159331 79598
rect 159633 79595 159699 79598
rect 161197 79595 161263 79598
rect 162526 79596 162532 79598
rect 162596 79596 162602 79660
rect 163078 79596 163084 79660
rect 163148 79658 163154 79660
rect 163589 79658 163655 79661
rect 163148 79656 163655 79658
rect 163148 79600 163594 79656
rect 163650 79600 163655 79656
rect 163148 79598 163655 79600
rect 163148 79596 163154 79598
rect 163589 79595 163655 79598
rect 164509 79656 164618 79661
rect 164509 79600 164514 79656
rect 164570 79600 164618 79656
rect 164509 79598 164618 79600
rect 164509 79595 164575 79598
rect 164918 79596 164924 79660
rect 164988 79658 164994 79660
rect 165478 79658 165538 79867
rect 167686 79661 167746 79901
rect 168046 79868 168052 79932
rect 168116 79930 168122 79932
rect 168327 79930 168332 79962
rect 168116 79906 168332 79930
rect 168388 79906 168393 79962
rect 170075 79962 170141 79967
rect 168695 79930 168761 79933
rect 169155 79932 169221 79933
rect 169150 79930 169156 79932
rect 168116 79901 168393 79906
rect 168560 79928 168761 79930
rect 168116 79870 168390 79901
rect 168560 79872 168700 79928
rect 168756 79872 168761 79928
rect 168560 79870 168761 79872
rect 169064 79870 169156 79930
rect 168116 79868 168122 79870
rect 168560 79794 168620 79870
rect 168695 79867 168761 79870
rect 169150 79868 169156 79870
rect 169220 79868 169226 79932
rect 169518 79868 169524 79932
rect 169588 79930 169594 79932
rect 169707 79930 169773 79933
rect 170075 79932 170080 79962
rect 170136 79932 170141 79962
rect 170351 79964 170417 79967
rect 170351 79962 170460 79964
rect 169588 79928 169773 79930
rect 169588 79872 169712 79928
rect 169768 79872 169773 79928
rect 169588 79870 169773 79872
rect 169588 79868 169594 79870
rect 169155 79867 169221 79868
rect 169707 79867 169773 79870
rect 170070 79868 170076 79932
rect 170140 79930 170146 79932
rect 170140 79870 170198 79930
rect 170351 79906 170356 79962
rect 170412 79906 170460 79962
rect 170995 79930 171061 79933
rect 170351 79901 170460 79906
rect 170140 79868 170146 79870
rect 170400 79797 170460 79901
rect 170630 79928 171061 79930
rect 170630 79872 171000 79928
rect 171056 79872 171061 79928
rect 170630 79870 171061 79872
rect 168741 79794 168807 79797
rect 168560 79792 168807 79794
rect 168560 79736 168746 79792
rect 168802 79736 168807 79792
rect 168560 79734 168807 79736
rect 168741 79731 168807 79734
rect 170397 79792 170463 79797
rect 170630 79796 170690 79870
rect 170995 79867 171061 79870
rect 171271 79930 171337 79933
rect 171412 79930 171472 80004
rect 171271 79928 171472 79930
rect 171271 79872 171276 79928
rect 171332 79872 171472 79928
rect 171731 79962 171797 79967
rect 171731 79906 171736 79962
rect 171792 79930 171797 79962
rect 173755 79962 173821 79967
rect 173387 79932 173453 79933
rect 173755 79932 173760 79962
rect 173816 79932 173821 79962
rect 174123 79962 174189 79967
rect 174123 79932 174128 79962
rect 174184 79932 174189 79962
rect 174675 79932 174741 79933
rect 172094 79930 172100 79932
rect 171792 79906 172100 79930
rect 171731 79901 172100 79906
rect 171271 79870 171472 79872
rect 171734 79870 172100 79901
rect 171271 79867 171337 79870
rect 172094 79868 172100 79870
rect 172164 79868 172170 79932
rect 173382 79930 173388 79932
rect 173296 79870 173388 79930
rect 173382 79868 173388 79870
rect 173452 79868 173458 79932
rect 173750 79868 173756 79932
rect 173820 79930 173826 79932
rect 173820 79870 173878 79930
rect 173820 79868 173826 79870
rect 174118 79868 174124 79932
rect 174188 79930 174194 79932
rect 174670 79930 174676 79932
rect 174188 79870 174246 79930
rect 174584 79870 174676 79930
rect 174188 79868 174194 79870
rect 174670 79868 174676 79870
rect 174740 79868 174746 79932
rect 174816 79930 174876 80006
rect 177024 80004 177068 80066
rect 177132 80004 177138 80068
rect 175227 79962 175293 79967
rect 174951 79930 175017 79933
rect 175227 79932 175232 79962
rect 175288 79932 175293 79962
rect 175411 79962 175477 79967
rect 174816 79928 175017 79930
rect 174816 79872 174956 79928
rect 175012 79872 175017 79928
rect 174816 79870 175017 79872
rect 173387 79867 173453 79868
rect 174675 79867 174741 79868
rect 174951 79867 175017 79870
rect 175222 79868 175228 79932
rect 175292 79930 175298 79932
rect 175292 79870 175350 79930
rect 175411 79906 175416 79962
rect 175472 79906 175477 79962
rect 175779 79962 175845 79967
rect 175779 79932 175784 79962
rect 175840 79932 175845 79962
rect 175411 79901 175477 79906
rect 175292 79868 175298 79870
rect 170397 79736 170402 79792
rect 170458 79736 170463 79792
rect 170397 79731 170463 79736
rect 170622 79732 170628 79796
rect 170692 79732 170698 79796
rect 171542 79732 171548 79796
rect 171612 79794 171618 79796
rect 172007 79794 172073 79797
rect 171612 79792 172073 79794
rect 171612 79736 172012 79792
rect 172068 79736 172073 79792
rect 171612 79734 172073 79736
rect 171612 79732 171618 79734
rect 172007 79731 172073 79734
rect 172513 79794 172579 79797
rect 174486 79794 174492 79796
rect 172513 79792 174492 79794
rect 172513 79736 172518 79792
rect 172574 79736 174492 79792
rect 172513 79734 174492 79736
rect 172513 79731 172579 79734
rect 174486 79732 174492 79734
rect 174556 79732 174562 79796
rect 174767 79794 174833 79797
rect 174905 79794 174971 79797
rect 174767 79792 174971 79794
rect 174767 79736 174772 79792
rect 174828 79736 174910 79792
rect 174966 79736 174971 79792
rect 174767 79734 174971 79736
rect 175414 79794 175474 79901
rect 175774 79868 175780 79932
rect 175844 79930 175850 79932
rect 176423 79930 176489 79933
rect 177024 79930 177084 80004
rect 179094 79967 179154 80142
rect 179091 79962 179157 79967
rect 177159 79930 177225 79933
rect 177987 79930 178053 79933
rect 178539 79932 178605 79933
rect 178534 79930 178540 79932
rect 175844 79870 175902 79930
rect 176423 79928 176946 79930
rect 176423 79872 176428 79928
rect 176484 79872 176946 79928
rect 176423 79870 176946 79872
rect 177024 79928 177225 79930
rect 177024 79872 177164 79928
rect 177220 79872 177225 79928
rect 177024 79870 177225 79872
rect 175844 79868 175850 79870
rect 176423 79867 176489 79870
rect 176326 79794 176332 79796
rect 175414 79734 176332 79794
rect 174767 79731 174833 79734
rect 174905 79731 174971 79734
rect 176326 79732 176332 79734
rect 176396 79732 176402 79796
rect 176886 79794 176946 79870
rect 177159 79867 177225 79870
rect 177806 79928 178053 79930
rect 177806 79872 177992 79928
rect 178048 79872 178053 79928
rect 177806 79870 178053 79872
rect 178448 79870 178540 79930
rect 177113 79794 177179 79797
rect 176886 79792 177179 79794
rect 176886 79736 177118 79792
rect 177174 79736 177179 79792
rect 176886 79734 177179 79736
rect 177113 79731 177179 79734
rect 164988 79598 165538 79658
rect 164988 79596 164994 79598
rect 166390 79596 166396 79660
rect 166460 79658 166466 79660
rect 166625 79658 166691 79661
rect 166460 79656 166691 79658
rect 166460 79600 166630 79656
rect 166686 79600 166691 79656
rect 166460 79598 166691 79600
rect 166460 79596 166466 79598
rect 166625 79595 166691 79598
rect 166758 79596 166764 79660
rect 166828 79658 166834 79660
rect 167361 79658 167427 79661
rect 166828 79656 167427 79658
rect 166828 79600 167366 79656
rect 167422 79600 167427 79656
rect 166828 79598 167427 79600
rect 166828 79596 166834 79598
rect 167361 79595 167427 79598
rect 167637 79656 167746 79661
rect 167637 79600 167642 79656
rect 167698 79600 167746 79656
rect 167637 79598 167746 79600
rect 167637 79595 167703 79598
rect 167862 79596 167868 79660
rect 167932 79658 167938 79660
rect 168097 79658 168163 79661
rect 177806 79658 177866 79870
rect 177987 79867 178053 79870
rect 178534 79868 178540 79870
rect 178604 79868 178610 79932
rect 179091 79906 179096 79962
rect 179152 79906 179157 79962
rect 179091 79901 179157 79906
rect 178539 79867 178605 79868
rect 177941 79794 178007 79797
rect 180609 79794 180675 79797
rect 177941 79792 180675 79794
rect 177941 79736 177946 79792
rect 178002 79736 180614 79792
rect 180670 79736 180675 79792
rect 177941 79734 180675 79736
rect 177941 79731 178007 79734
rect 180609 79731 180675 79734
rect 178033 79660 178099 79661
rect 167932 79656 168163 79658
rect 167932 79600 168102 79656
rect 168158 79600 168163 79656
rect 167932 79598 168163 79600
rect 167932 79596 167938 79598
rect 168097 79595 168163 79598
rect 168330 79598 177866 79658
rect 71773 79522 71839 79525
rect 168330 79522 168390 79598
rect 177982 79596 177988 79660
rect 178052 79658 178099 79660
rect 178052 79656 178144 79658
rect 178094 79600 178144 79656
rect 178052 79598 178144 79600
rect 178052 79596 178099 79598
rect 178033 79595 178099 79596
rect 168557 79524 168623 79525
rect 170489 79524 170555 79525
rect 168557 79522 168604 79524
rect 71773 79520 168390 79522
rect 71773 79464 71778 79520
rect 71834 79464 168390 79520
rect 71773 79462 168390 79464
rect 168512 79520 168604 79522
rect 168512 79464 168562 79520
rect 168512 79462 168604 79464
rect 71773 79459 71839 79462
rect 168557 79460 168604 79462
rect 168668 79460 168674 79524
rect 170438 79522 170444 79524
rect 170398 79462 170444 79522
rect 170508 79520 170555 79524
rect 170550 79464 170555 79520
rect 170438 79460 170444 79462
rect 170508 79460 170555 79464
rect 171910 79460 171916 79524
rect 171980 79522 171986 79524
rect 172421 79522 172487 79525
rect 173341 79524 173407 79525
rect 173341 79522 173388 79524
rect 171980 79520 172487 79522
rect 171980 79464 172426 79520
rect 172482 79464 172487 79520
rect 171980 79462 172487 79464
rect 173296 79520 173388 79522
rect 173296 79464 173346 79520
rect 173296 79462 173388 79464
rect 171980 79460 171986 79462
rect 168557 79459 168623 79460
rect 170489 79459 170555 79460
rect 172421 79459 172487 79462
rect 173341 79460 173388 79462
rect 173452 79460 173458 79524
rect 177665 79522 177731 79525
rect 331213 79522 331279 79525
rect 177665 79520 331279 79522
rect 177665 79464 177670 79520
rect 177726 79464 331218 79520
rect 331274 79464 331279 79520
rect 177665 79462 331279 79464
rect 173341 79459 173407 79460
rect 177665 79459 177731 79462
rect 331213 79459 331279 79462
rect 116577 79386 116643 79389
rect 177205 79386 177271 79389
rect 580206 79386 580212 79388
rect 116577 79384 176026 79386
rect 116577 79328 116582 79384
rect 116638 79328 176026 79384
rect 116577 79326 176026 79328
rect 116577 79323 116643 79326
rect 3417 79250 3483 79253
rect 175966 79250 176026 79326
rect 177205 79384 580212 79386
rect 177205 79328 177210 79384
rect 177266 79328 580212 79384
rect 177205 79326 580212 79328
rect 177205 79323 177271 79326
rect 580206 79324 580212 79326
rect 580276 79324 580282 79388
rect 178217 79250 178283 79253
rect 3417 79248 175888 79250
rect 3417 79192 3422 79248
rect 3478 79192 175888 79248
rect 3417 79190 175888 79192
rect 175966 79248 178283 79250
rect 175966 79192 178222 79248
rect 178278 79192 178283 79248
rect 175966 79190 178283 79192
rect 3417 79187 3483 79190
rect 135897 79114 135963 79117
rect 149237 79114 149303 79117
rect 135897 79112 149303 79114
rect 135897 79056 135902 79112
rect 135958 79056 149242 79112
rect 149298 79056 149303 79112
rect 135897 79054 149303 79056
rect 135897 79051 135963 79054
rect 149237 79051 149303 79054
rect 155534 79052 155540 79116
rect 155604 79114 155610 79116
rect 157425 79114 157491 79117
rect 155604 79112 157491 79114
rect 155604 79056 157430 79112
rect 157486 79056 157491 79112
rect 155604 79054 157491 79056
rect 155604 79052 155610 79054
rect 157425 79051 157491 79054
rect 162158 79052 162164 79116
rect 162228 79114 162234 79116
rect 162853 79114 162919 79117
rect 162228 79112 162919 79114
rect 162228 79056 162858 79112
rect 162914 79056 162919 79112
rect 162228 79054 162919 79056
rect 162228 79052 162234 79054
rect 162853 79051 162919 79054
rect 163497 79114 163563 79117
rect 163630 79114 163636 79116
rect 163497 79112 163636 79114
rect 163497 79056 163502 79112
rect 163558 79056 163636 79112
rect 163497 79054 163636 79056
rect 163497 79051 163563 79054
rect 163630 79052 163636 79054
rect 163700 79052 163706 79116
rect 165613 79114 165679 79117
rect 168097 79114 168163 79117
rect 165613 79112 168163 79114
rect 165613 79056 165618 79112
rect 165674 79056 168102 79112
rect 168158 79056 168163 79112
rect 165613 79054 168163 79056
rect 165613 79051 165679 79054
rect 168097 79051 168163 79054
rect 168557 79114 168623 79117
rect 168557 79112 173910 79114
rect 168557 79056 168562 79112
rect 168618 79056 173910 79112
rect 168557 79054 173910 79056
rect 168557 79051 168623 79054
rect 138197 78978 138263 78981
rect 156689 78980 156755 78981
rect 138974 78978 138980 78980
rect 138197 78976 138980 78978
rect 138197 78920 138202 78976
rect 138258 78920 138980 78976
rect 138197 78918 138980 78920
rect 138197 78915 138263 78918
rect 138974 78916 138980 78918
rect 139044 78916 139050 78980
rect 156638 78916 156644 78980
rect 156708 78978 156755 78980
rect 158621 78978 158687 78981
rect 162301 78980 162367 78981
rect 164049 78980 164115 78981
rect 158846 78978 158852 78980
rect 156708 78976 156800 78978
rect 156750 78920 156800 78976
rect 156708 78918 156800 78920
rect 158621 78976 158852 78978
rect 158621 78920 158626 78976
rect 158682 78920 158852 78976
rect 158621 78918 158852 78920
rect 156708 78916 156755 78918
rect 156689 78915 156755 78916
rect 158621 78915 158687 78918
rect 158846 78916 158852 78918
rect 158916 78916 158922 78980
rect 162301 78978 162348 78980
rect 162256 78976 162348 78978
rect 162256 78920 162306 78976
rect 162256 78918 162348 78920
rect 162301 78916 162348 78918
rect 162412 78916 162418 78980
rect 163998 78916 164004 78980
rect 164068 78978 164115 78980
rect 164417 78978 164483 78981
rect 164068 78976 164160 78978
rect 164110 78920 164160 78976
rect 164068 78918 164160 78920
rect 164417 78976 167010 78978
rect 164417 78920 164422 78976
rect 164478 78920 167010 78976
rect 164417 78918 167010 78920
rect 164068 78916 164115 78918
rect 162301 78915 162367 78916
rect 164049 78915 164115 78916
rect 164417 78915 164483 78918
rect 136265 78842 136331 78845
rect 134566 78840 136331 78842
rect 134566 78784 136270 78840
rect 136326 78784 136331 78840
rect 134566 78782 136331 78784
rect 133965 78706 134031 78709
rect 134566 78706 134626 78782
rect 136265 78779 136331 78782
rect 136582 78780 136588 78844
rect 136652 78842 136658 78844
rect 137737 78842 137803 78845
rect 136652 78840 137803 78842
rect 136652 78784 137742 78840
rect 137798 78784 137803 78840
rect 136652 78782 137803 78784
rect 136652 78780 136658 78782
rect 137737 78779 137803 78782
rect 138054 78780 138060 78844
rect 138124 78842 138130 78844
rect 138381 78842 138447 78845
rect 138124 78840 138447 78842
rect 138124 78784 138386 78840
rect 138442 78784 138447 78840
rect 138124 78782 138447 78784
rect 138124 78780 138130 78782
rect 138381 78779 138447 78782
rect 160686 78780 160692 78844
rect 160756 78842 160762 78844
rect 161105 78842 161171 78845
rect 161565 78842 161631 78845
rect 161933 78844 161999 78845
rect 161933 78842 161980 78844
rect 160756 78840 161171 78842
rect 160756 78784 161110 78840
rect 161166 78784 161171 78840
rect 160756 78782 161171 78784
rect 160756 78780 160762 78782
rect 161105 78779 161171 78782
rect 161430 78840 161631 78842
rect 161430 78784 161570 78840
rect 161626 78784 161631 78840
rect 161430 78782 161631 78784
rect 161888 78840 161980 78842
rect 161888 78784 161938 78840
rect 161888 78782 161980 78784
rect 133965 78704 134626 78706
rect 133965 78648 133970 78704
rect 134026 78648 134626 78704
rect 133965 78646 134626 78648
rect 133965 78643 134031 78646
rect 134926 78644 134932 78708
rect 134996 78706 135002 78708
rect 135069 78706 135135 78709
rect 136173 78708 136239 78709
rect 136173 78706 136220 78708
rect 134996 78704 135135 78706
rect 134996 78648 135074 78704
rect 135130 78648 135135 78704
rect 134996 78646 135135 78648
rect 136128 78704 136220 78706
rect 136128 78648 136178 78704
rect 136128 78646 136220 78648
rect 134996 78644 135002 78646
rect 135069 78643 135135 78646
rect 136173 78644 136220 78646
rect 136284 78644 136290 78708
rect 136725 78706 136791 78709
rect 137737 78708 137803 78709
rect 137502 78706 137508 78708
rect 136725 78704 137508 78706
rect 136725 78648 136730 78704
rect 136786 78648 137508 78704
rect 136725 78646 137508 78648
rect 136173 78643 136239 78644
rect 136725 78643 136791 78646
rect 137502 78644 137508 78646
rect 137572 78644 137578 78708
rect 137686 78644 137692 78708
rect 137756 78706 137803 78708
rect 138105 78706 138171 78709
rect 139485 78708 139551 78709
rect 138238 78706 138244 78708
rect 137756 78704 137848 78706
rect 137798 78648 137848 78704
rect 137756 78646 137848 78648
rect 138105 78704 138244 78706
rect 138105 78648 138110 78704
rect 138166 78648 138244 78704
rect 138105 78646 138244 78648
rect 137756 78644 137803 78646
rect 137737 78643 137803 78644
rect 138105 78643 138171 78646
rect 138238 78644 138244 78646
rect 138308 78644 138314 78708
rect 139485 78704 139532 78708
rect 139596 78706 139602 78708
rect 141233 78706 141299 78709
rect 141366 78706 141372 78708
rect 139485 78648 139490 78704
rect 139485 78644 139532 78648
rect 139596 78646 139642 78706
rect 141233 78704 141372 78706
rect 141233 78648 141238 78704
rect 141294 78648 141372 78704
rect 141233 78646 141372 78648
rect 139596 78644 139602 78646
rect 139485 78643 139551 78644
rect 141233 78643 141299 78646
rect 141366 78644 141372 78646
rect 141436 78644 141442 78708
rect 160870 78644 160876 78708
rect 160940 78706 160946 78708
rect 161430 78706 161490 78782
rect 161565 78779 161631 78782
rect 161933 78780 161980 78782
rect 162044 78780 162050 78844
rect 163262 78780 163268 78844
rect 163332 78842 163338 78844
rect 164141 78842 164207 78845
rect 163332 78840 164207 78842
rect 163332 78784 164146 78840
rect 164202 78784 164207 78840
rect 163332 78782 164207 78784
rect 163332 78780 163338 78782
rect 161933 78779 161999 78780
rect 164141 78779 164207 78782
rect 166441 78842 166507 78845
rect 166717 78844 166783 78845
rect 166574 78842 166580 78844
rect 166441 78840 166580 78842
rect 166441 78784 166446 78840
rect 166502 78784 166580 78840
rect 166441 78782 166580 78784
rect 166441 78779 166507 78782
rect 166574 78780 166580 78782
rect 166644 78780 166650 78844
rect 166717 78840 166764 78844
rect 166828 78842 166834 78844
rect 166950 78842 167010 78918
rect 167678 78916 167684 78980
rect 167748 78978 167754 78980
rect 168281 78978 168347 78981
rect 167748 78976 168347 78978
rect 167748 78920 168286 78976
rect 168342 78920 168347 78976
rect 167748 78918 168347 78920
rect 173850 78978 173910 79054
rect 174854 79052 174860 79116
rect 174924 79114 174930 79116
rect 175181 79114 175247 79117
rect 174924 79112 175247 79114
rect 174924 79056 175186 79112
rect 175242 79056 175247 79112
rect 174924 79054 175247 79056
rect 175828 79114 175888 79190
rect 178217 79187 178283 79190
rect 178401 79250 178467 79253
rect 178534 79250 178540 79252
rect 178401 79248 178540 79250
rect 178401 79192 178406 79248
rect 178462 79192 178540 79248
rect 178401 79190 178540 79192
rect 178401 79187 178467 79190
rect 178534 79188 178540 79190
rect 178604 79188 178610 79252
rect 177113 79114 177179 79117
rect 175828 79112 177179 79114
rect 175828 79056 177118 79112
rect 177174 79056 177179 79112
rect 175828 79054 177179 79056
rect 174924 79052 174930 79054
rect 175181 79051 175247 79054
rect 177113 79051 177179 79054
rect 177481 79114 177547 79117
rect 397453 79114 397519 79117
rect 177481 79112 397519 79114
rect 177481 79056 177486 79112
rect 177542 79056 397458 79112
rect 397514 79056 397519 79112
rect 177481 79054 397519 79056
rect 177481 79051 177547 79054
rect 397453 79051 397519 79054
rect 178493 78978 178559 78981
rect 173850 78976 178559 78978
rect 173850 78920 178498 78976
rect 178554 78920 178559 78976
rect 173850 78918 178559 78920
rect 167748 78916 167754 78918
rect 168281 78915 168347 78918
rect 178493 78915 178559 78918
rect 180517 78978 180583 78981
rect 462313 78978 462379 78981
rect 180517 78976 462379 78978
rect 180517 78920 180522 78976
rect 180578 78920 462318 78976
rect 462374 78920 462379 78976
rect 180517 78918 462379 78920
rect 180517 78915 180583 78918
rect 462313 78915 462379 78918
rect 176653 78842 176719 78845
rect 166717 78784 166722 78840
rect 166717 78780 166764 78784
rect 166828 78782 166874 78842
rect 166950 78840 176719 78842
rect 166950 78784 176658 78840
rect 176714 78784 176719 78840
rect 166950 78782 176719 78784
rect 166828 78780 166834 78782
rect 166717 78779 166783 78780
rect 176653 78779 176719 78782
rect 176929 78842 176995 78845
rect 580533 78842 580599 78845
rect 176929 78840 580599 78842
rect 176929 78784 176934 78840
rect 176990 78784 580538 78840
rect 580594 78784 580599 78840
rect 176929 78782 580599 78784
rect 176929 78779 176995 78782
rect 580533 78779 580599 78782
rect 160940 78646 161490 78706
rect 160940 78644 160946 78646
rect 161606 78644 161612 78708
rect 161676 78706 161682 78708
rect 161841 78706 161907 78709
rect 161676 78704 161907 78706
rect 161676 78648 161846 78704
rect 161902 78648 161907 78704
rect 161676 78646 161907 78648
rect 161676 78644 161682 78646
rect 161841 78643 161907 78646
rect 162342 78644 162348 78708
rect 162412 78706 162418 78708
rect 162485 78706 162551 78709
rect 162412 78704 162551 78706
rect 162412 78648 162490 78704
rect 162546 78648 162551 78704
rect 162412 78646 162551 78648
rect 162412 78644 162418 78646
rect 162485 78643 162551 78646
rect 163078 78644 163084 78708
rect 163148 78706 163154 78708
rect 163313 78706 163379 78709
rect 163148 78704 163379 78706
rect 163148 78648 163318 78704
rect 163374 78648 163379 78704
rect 163148 78646 163379 78648
rect 163148 78644 163154 78646
rect 163313 78643 163379 78646
rect 163446 78644 163452 78708
rect 163516 78706 163522 78708
rect 163957 78706 164023 78709
rect 163516 78704 164023 78706
rect 163516 78648 163962 78704
rect 164018 78648 164023 78704
rect 163516 78646 164023 78648
rect 163516 78644 163522 78646
rect 163957 78643 164023 78646
rect 165102 78644 165108 78708
rect 165172 78706 165178 78708
rect 165245 78706 165311 78709
rect 165521 78708 165587 78709
rect 165470 78706 165476 78708
rect 165172 78704 165311 78706
rect 165172 78648 165250 78704
rect 165306 78648 165311 78704
rect 165172 78646 165311 78648
rect 165430 78646 165476 78706
rect 165540 78704 165587 78708
rect 165582 78648 165587 78704
rect 165172 78644 165178 78646
rect 165245 78643 165311 78646
rect 165470 78644 165476 78646
rect 165540 78644 165587 78648
rect 166574 78644 166580 78708
rect 166644 78706 166650 78708
rect 166901 78706 166967 78709
rect 166644 78704 166967 78706
rect 166644 78648 166906 78704
rect 166962 78648 166967 78704
rect 166644 78646 166967 78648
rect 166644 78644 166650 78646
rect 165521 78643 165587 78644
rect 166901 78643 166967 78646
rect 167494 78644 167500 78708
rect 167564 78706 167570 78708
rect 168189 78706 168255 78709
rect 167564 78704 168255 78706
rect 167564 78648 168194 78704
rect 168250 78648 168255 78704
rect 167564 78646 168255 78648
rect 167564 78644 167570 78646
rect 168189 78643 168255 78646
rect 169661 78708 169727 78709
rect 171041 78708 171107 78709
rect 169661 78704 169708 78708
rect 169772 78706 169778 78708
rect 170990 78706 170996 78708
rect 169661 78648 169666 78704
rect 169661 78644 169708 78648
rect 169772 78646 169818 78706
rect 170950 78646 170996 78706
rect 171060 78704 171107 78708
rect 171102 78648 171107 78704
rect 169772 78644 169778 78646
rect 170990 78644 170996 78646
rect 171060 78644 171107 78648
rect 171726 78644 171732 78708
rect 171796 78706 171802 78708
rect 172145 78706 172211 78709
rect 175181 78708 175247 78709
rect 176009 78708 176075 78709
rect 175181 78706 175228 78708
rect 171796 78704 172211 78706
rect 171796 78648 172150 78704
rect 172206 78648 172211 78704
rect 171796 78646 172211 78648
rect 175136 78704 175228 78706
rect 175136 78648 175186 78704
rect 175136 78646 175228 78648
rect 171796 78644 171802 78646
rect 169661 78643 169727 78644
rect 171041 78643 171107 78644
rect 172145 78643 172211 78646
rect 175181 78644 175228 78646
rect 175292 78644 175298 78708
rect 175958 78706 175964 78708
rect 175918 78646 175964 78706
rect 176028 78704 176075 78708
rect 176070 78648 176075 78704
rect 175958 78644 175964 78646
rect 176028 78644 176075 78648
rect 175181 78643 175247 78644
rect 176009 78643 176075 78644
rect 176561 78706 176627 78709
rect 580717 78706 580783 78709
rect 176561 78704 580783 78706
rect 176561 78648 176566 78704
rect 176622 78648 580722 78704
rect 580778 78648 580783 78704
rect 176561 78646 580783 78648
rect 176561 78643 176627 78646
rect 580717 78643 580783 78646
rect 4061 78570 4127 78573
rect 172145 78572 172211 78573
rect 4061 78568 171610 78570
rect 4061 78512 4066 78568
rect 4122 78512 171610 78568
rect 4061 78510 171610 78512
rect 4061 78507 4127 78510
rect 119337 78434 119403 78437
rect 170949 78434 171015 78437
rect 119337 78432 171015 78434
rect 119337 78376 119342 78432
rect 119398 78376 170954 78432
rect 171010 78376 171015 78432
rect 119337 78374 171015 78376
rect 119337 78371 119403 78374
rect 170949 78371 171015 78374
rect 150750 78236 150756 78300
rect 150820 78298 150826 78300
rect 150985 78298 151051 78301
rect 150820 78296 151051 78298
rect 150820 78240 150990 78296
rect 151046 78240 151051 78296
rect 150820 78238 151051 78240
rect 150820 78236 150826 78238
rect 150985 78235 151051 78238
rect 166206 78236 166212 78300
rect 166276 78298 166282 78300
rect 166809 78298 166875 78301
rect 166276 78296 166875 78298
rect 166276 78240 166814 78296
rect 166870 78240 166875 78296
rect 166276 78238 166875 78240
rect 171550 78298 171610 78510
rect 172094 78508 172100 78572
rect 172164 78570 172211 78572
rect 174169 78570 174235 78573
rect 179873 78570 179939 78573
rect 172164 78568 172256 78570
rect 172206 78512 172256 78568
rect 172164 78510 172256 78512
rect 174169 78568 179939 78570
rect 174169 78512 174174 78568
rect 174230 78512 179878 78568
rect 179934 78512 179939 78568
rect 174169 78510 179939 78512
rect 172164 78508 172211 78510
rect 172145 78507 172211 78508
rect 174169 78507 174235 78510
rect 179873 78507 179939 78510
rect 172094 78372 172100 78436
rect 172164 78434 172170 78436
rect 172329 78434 172395 78437
rect 172164 78432 172395 78434
rect 172164 78376 172334 78432
rect 172390 78376 172395 78432
rect 172164 78374 172395 78376
rect 172164 78372 172170 78374
rect 172329 78371 172395 78374
rect 174261 78434 174327 78437
rect 174670 78434 174676 78436
rect 174261 78432 174676 78434
rect 174261 78376 174266 78432
rect 174322 78376 174676 78432
rect 174261 78374 174676 78376
rect 174261 78371 174327 78374
rect 174670 78372 174676 78374
rect 174740 78372 174746 78436
rect 175549 78434 175615 78437
rect 176510 78434 176516 78436
rect 175549 78432 176516 78434
rect 175549 78376 175554 78432
rect 175610 78376 176516 78432
rect 175549 78374 176516 78376
rect 175549 78371 175615 78374
rect 176510 78372 176516 78374
rect 176580 78372 176586 78436
rect 179689 78434 179755 78437
rect 176886 78432 179755 78434
rect 176886 78376 179694 78432
rect 179750 78376 179755 78432
rect 176886 78374 179755 78376
rect 176886 78298 176946 78374
rect 179689 78371 179755 78374
rect 171550 78238 176946 78298
rect 177021 78298 177087 78301
rect 188981 78298 189047 78301
rect 177021 78296 189047 78298
rect 177021 78240 177026 78296
rect 177082 78240 188986 78296
rect 189042 78240 189047 78296
rect 177021 78238 189047 78240
rect 166276 78236 166282 78238
rect 166809 78235 166875 78238
rect 177021 78235 177087 78238
rect 188981 78235 189047 78238
rect 131389 78162 131455 78165
rect 132861 78164 132927 78165
rect 132350 78162 132356 78164
rect 131389 78160 132356 78162
rect 131389 78104 131394 78160
rect 131450 78104 132356 78160
rect 131389 78102 132356 78104
rect 131389 78099 131455 78102
rect 132350 78100 132356 78102
rect 132420 78100 132426 78164
rect 132861 78162 132908 78164
rect 132816 78160 132908 78162
rect 132816 78104 132866 78160
rect 132816 78102 132908 78104
rect 132861 78100 132908 78102
rect 132972 78100 132978 78164
rect 139158 78100 139164 78164
rect 139228 78162 139234 78164
rect 151261 78162 151327 78165
rect 139228 78160 151327 78162
rect 139228 78104 151266 78160
rect 151322 78104 151327 78160
rect 139228 78102 151327 78104
rect 139228 78100 139234 78102
rect 132861 78099 132927 78100
rect 151261 78099 151327 78102
rect 167310 78100 167316 78164
rect 167380 78162 167386 78164
rect 167545 78162 167611 78165
rect 167380 78160 167611 78162
rect 167380 78104 167550 78160
rect 167606 78104 167611 78160
rect 167380 78102 167611 78104
rect 167380 78100 167386 78102
rect 167545 78099 167611 78102
rect 174302 78100 174308 78164
rect 174372 78162 174378 78164
rect 174670 78162 174676 78164
rect 174372 78102 174676 78162
rect 174372 78100 174378 78102
rect 174670 78100 174676 78102
rect 174740 78100 174746 78164
rect 177113 78162 177179 78165
rect 178309 78162 178375 78165
rect 177113 78160 178375 78162
rect 177113 78104 177118 78160
rect 177174 78104 178314 78160
rect 178370 78104 178375 78160
rect 177113 78102 178375 78104
rect 177113 78099 177179 78102
rect 178309 78099 178375 78102
rect 124857 78026 124923 78029
rect 133321 78026 133387 78029
rect 124857 78024 133387 78026
rect 124857 77968 124862 78024
rect 124918 77968 133326 78024
rect 133382 77968 133387 78024
rect 124857 77966 133387 77968
rect 124857 77963 124923 77966
rect 133321 77963 133387 77966
rect 165429 78026 165495 78029
rect 178033 78026 178099 78029
rect 165429 78024 178099 78026
rect 165429 77968 165434 78024
rect 165490 77968 178038 78024
rect 178094 77968 178099 78024
rect 165429 77966 178099 77968
rect 165429 77963 165495 77966
rect 178033 77963 178099 77966
rect 95877 77890 95943 77893
rect 131982 77890 131988 77892
rect 95877 77888 131988 77890
rect 95877 77832 95882 77888
rect 95938 77832 131988 77888
rect 95877 77830 131988 77832
rect 95877 77827 95943 77830
rect 131982 77828 131988 77830
rect 132052 77828 132058 77892
rect 136725 77890 136791 77893
rect 137870 77890 137876 77892
rect 136725 77888 137876 77890
rect 136725 77832 136730 77888
rect 136786 77832 137876 77888
rect 136725 77830 137876 77832
rect 136725 77827 136791 77830
rect 137870 77828 137876 77830
rect 137940 77828 137946 77892
rect 170254 77828 170260 77892
rect 170324 77890 170330 77892
rect 170673 77890 170739 77893
rect 174169 77892 174235 77893
rect 170324 77888 170739 77890
rect 170324 77832 170678 77888
rect 170734 77832 170739 77888
rect 170324 77830 170739 77832
rect 170324 77828 170330 77830
rect 170673 77827 170739 77830
rect 174118 77828 174124 77892
rect 174188 77890 174235 77892
rect 174629 77890 174695 77893
rect 176878 77890 176884 77892
rect 174188 77888 174280 77890
rect 174230 77832 174280 77888
rect 174188 77830 174280 77832
rect 174629 77888 176884 77890
rect 174629 77832 174634 77888
rect 174690 77832 176884 77888
rect 174629 77830 176884 77832
rect 174188 77828 174235 77830
rect 174169 77827 174235 77828
rect 174629 77827 174695 77830
rect 176878 77828 176884 77830
rect 176948 77828 176954 77892
rect 129641 77754 129707 77757
rect 154389 77754 154455 77757
rect 129641 77752 154455 77754
rect 129641 77696 129646 77752
rect 129702 77696 154394 77752
rect 154450 77696 154455 77752
rect 129641 77694 154455 77696
rect 129641 77691 129707 77694
rect 154389 77691 154455 77694
rect 170949 77754 171015 77757
rect 176469 77754 176535 77757
rect 177573 77754 177639 77757
rect 170949 77752 176535 77754
rect 170949 77696 170954 77752
rect 171010 77696 176474 77752
rect 176530 77696 176535 77752
rect 170949 77694 176535 77696
rect 170949 77691 171015 77694
rect 176469 77691 176535 77694
rect 176610 77752 177639 77754
rect 176610 77696 177578 77752
rect 177634 77696 177639 77752
rect 176610 77694 177639 77696
rect 140865 77618 140931 77621
rect 140998 77618 141004 77620
rect 140865 77616 141004 77618
rect 140865 77560 140870 77616
rect 140926 77560 141004 77616
rect 140865 77558 141004 77560
rect 140865 77555 140931 77558
rect 140998 77556 141004 77558
rect 141068 77556 141074 77620
rect 144085 77618 144151 77621
rect 144494 77618 144500 77620
rect 144085 77616 144500 77618
rect 144085 77560 144090 77616
rect 144146 77560 144500 77616
rect 144085 77558 144500 77560
rect 144085 77555 144151 77558
rect 144494 77556 144500 77558
rect 144564 77556 144570 77620
rect 168005 77618 168071 77621
rect 176610 77618 176670 77694
rect 177573 77691 177639 77694
rect 168005 77616 174002 77618
rect 168005 77560 168010 77616
rect 168066 77560 174002 77616
rect 168005 77558 174002 77560
rect 168005 77555 168071 77558
rect 142838 77420 142844 77484
rect 142908 77482 142914 77484
rect 143349 77482 143415 77485
rect 142908 77480 143415 77482
rect 142908 77424 143354 77480
rect 143410 77424 143415 77480
rect 142908 77422 143415 77424
rect 142908 77420 142914 77422
rect 143349 77419 143415 77422
rect 144310 77420 144316 77484
rect 144380 77482 144386 77484
rect 144545 77482 144611 77485
rect 144380 77480 144611 77482
rect 144380 77424 144550 77480
rect 144606 77424 144611 77480
rect 144380 77422 144611 77424
rect 144380 77420 144386 77422
rect 144545 77419 144611 77422
rect 144913 77482 144979 77485
rect 145230 77482 145236 77484
rect 144913 77480 145236 77482
rect 144913 77424 144918 77480
rect 144974 77424 145236 77480
rect 144913 77422 145236 77424
rect 144913 77419 144979 77422
rect 145230 77420 145236 77422
rect 145300 77420 145306 77484
rect 145414 77420 145420 77484
rect 145484 77482 145490 77484
rect 145649 77482 145715 77485
rect 146201 77482 146267 77485
rect 147489 77484 147555 77485
rect 147438 77482 147444 77484
rect 145484 77480 145715 77482
rect 145484 77424 145654 77480
rect 145710 77424 145715 77480
rect 145484 77422 145715 77424
rect 145484 77420 145490 77422
rect 145649 77419 145715 77422
rect 145790 77480 146267 77482
rect 145790 77424 146206 77480
rect 146262 77424 146267 77480
rect 145790 77422 146267 77424
rect 147398 77422 147444 77482
rect 147508 77480 147555 77484
rect 147550 77424 147555 77480
rect 135529 77348 135595 77349
rect 135478 77284 135484 77348
rect 135548 77346 135595 77348
rect 135548 77344 135640 77346
rect 135590 77288 135640 77344
rect 135548 77286 135640 77288
rect 135548 77284 135595 77286
rect 140630 77284 140636 77348
rect 140700 77346 140706 77348
rect 140700 77286 142906 77346
rect 140700 77284 140706 77286
rect 135529 77283 135595 77284
rect 131021 77210 131087 77213
rect 131614 77210 131620 77212
rect 131021 77208 131620 77210
rect 131021 77152 131026 77208
rect 131082 77152 131620 77208
rect 131021 77150 131620 77152
rect 131021 77147 131087 77150
rect 131614 77148 131620 77150
rect 131684 77148 131690 77212
rect 142846 77210 142906 77286
rect 143022 77284 143028 77348
rect 143092 77346 143098 77348
rect 143257 77346 143323 77349
rect 143092 77344 143323 77346
rect 143092 77288 143262 77344
rect 143318 77288 143323 77344
rect 143092 77286 143323 77288
rect 143092 77284 143098 77286
rect 143257 77283 143323 77286
rect 145230 77284 145236 77348
rect 145300 77346 145306 77348
rect 145790 77346 145850 77422
rect 146201 77419 146267 77422
rect 147438 77420 147444 77422
rect 147508 77420 147555 77424
rect 147489 77419 147555 77420
rect 145300 77286 145850 77346
rect 146569 77346 146635 77349
rect 146886 77346 146892 77348
rect 146569 77344 146892 77346
rect 146569 77288 146574 77344
rect 146630 77288 146892 77344
rect 146569 77286 146892 77288
rect 145300 77284 145306 77286
rect 146569 77283 146635 77286
rect 146886 77284 146892 77286
rect 146956 77284 146962 77348
rect 147254 77284 147260 77348
rect 147324 77346 147330 77348
rect 147397 77346 147463 77349
rect 161289 77348 161355 77349
rect 161238 77346 161244 77348
rect 147324 77344 147463 77346
rect 147324 77288 147402 77344
rect 147458 77288 147463 77344
rect 147324 77286 147463 77288
rect 161198 77286 161244 77346
rect 161308 77344 161355 77348
rect 161350 77288 161355 77344
rect 147324 77284 147330 77286
rect 147397 77283 147463 77286
rect 161238 77284 161244 77286
rect 161308 77284 161355 77288
rect 173566 77284 173572 77348
rect 173636 77346 173642 77348
rect 173709 77346 173775 77349
rect 173636 77344 173775 77346
rect 173636 77288 173714 77344
rect 173770 77288 173775 77344
rect 173636 77286 173775 77288
rect 173942 77346 174002 77558
rect 176150 77558 176670 77618
rect 176150 77482 176210 77558
rect 177062 77556 177068 77620
rect 177132 77618 177138 77620
rect 189349 77618 189415 77621
rect 177132 77616 189415 77618
rect 177132 77560 189354 77616
rect 189410 77560 189415 77616
rect 177132 77558 189415 77560
rect 177132 77556 177138 77558
rect 189349 77555 189415 77558
rect 175230 77422 176210 77482
rect 176469 77482 176535 77485
rect 179045 77482 179111 77485
rect 176469 77480 179111 77482
rect 176469 77424 176474 77480
rect 176530 77424 179050 77480
rect 179106 77424 179111 77480
rect 176469 77422 179111 77424
rect 173942 77286 174738 77346
rect 173636 77284 173642 77286
rect 161289 77283 161355 77284
rect 173709 77283 173775 77286
rect 152181 77210 152247 77213
rect 170397 77212 170463 77213
rect 170397 77210 170444 77212
rect 142846 77208 152247 77210
rect 142846 77152 152186 77208
rect 152242 77152 152247 77208
rect 142846 77150 152247 77152
rect 170352 77208 170444 77210
rect 170352 77152 170402 77208
rect 170352 77150 170444 77152
rect 152181 77147 152247 77150
rect 170397 77148 170444 77150
rect 170508 77148 170514 77212
rect 174678 77210 174738 77286
rect 175230 77210 175290 77422
rect 176469 77419 176535 77422
rect 179045 77419 179111 77422
rect 176837 77346 176903 77349
rect 189073 77346 189139 77349
rect 176837 77344 189139 77346
rect 176837 77288 176842 77344
rect 176898 77288 189078 77344
rect 189134 77288 189139 77344
rect 176837 77286 189139 77288
rect 176837 77283 176903 77286
rect 189073 77283 189139 77286
rect 174678 77150 175290 77210
rect 170397 77147 170463 77148
rect 153745 77074 153811 77077
rect 153878 77074 153884 77076
rect 153745 77072 153884 77074
rect 153745 77016 153750 77072
rect 153806 77016 153884 77072
rect 153745 77014 153884 77016
rect 153745 77011 153811 77014
rect 153878 77012 153884 77014
rect 153948 77012 153954 77076
rect 154297 77074 154363 77077
rect 303613 77074 303679 77077
rect 154297 77072 303679 77074
rect 154297 77016 154302 77072
rect 154358 77016 303618 77072
rect 303674 77016 303679 77072
rect 154297 77014 303679 77016
rect 154297 77011 154363 77014
rect 303613 77011 303679 77014
rect 157926 76876 157932 76940
rect 157996 76938 158002 76940
rect 158437 76938 158503 76941
rect 157996 76936 158503 76938
rect 157996 76880 158442 76936
rect 158498 76880 158503 76936
rect 157996 76878 158503 76880
rect 157996 76876 158002 76878
rect 158437 76875 158503 76878
rect 160093 76938 160159 76941
rect 160502 76938 160508 76940
rect 160093 76936 160508 76938
rect 160093 76880 160098 76936
rect 160154 76880 160508 76936
rect 160093 76878 160508 76880
rect 160093 76875 160159 76878
rect 160502 76876 160508 76878
rect 160572 76876 160578 76940
rect 163589 76938 163655 76941
rect 419533 76938 419599 76941
rect 163589 76936 419599 76938
rect 163589 76880 163594 76936
rect 163650 76880 419538 76936
rect 419594 76880 419599 76936
rect 163589 76878 419599 76880
rect 163589 76875 163655 76878
rect 419533 76875 419599 76878
rect 145598 76740 145604 76804
rect 145668 76802 145674 76804
rect 149421 76802 149487 76805
rect 145668 76800 149487 76802
rect 145668 76744 149426 76800
rect 149482 76744 149487 76800
rect 145668 76742 149487 76744
rect 145668 76740 145674 76742
rect 149421 76739 149487 76742
rect 176285 76802 176351 76805
rect 451273 76802 451339 76805
rect 176285 76800 451339 76802
rect 176285 76744 176290 76800
rect 176346 76744 451278 76800
rect 451334 76744 451339 76800
rect 176285 76742 451339 76744
rect 176285 76739 176351 76742
rect 451273 76739 451339 76742
rect 140998 76604 141004 76668
rect 141068 76666 141074 76668
rect 142061 76666 142127 76669
rect 141068 76664 142127 76666
rect 141068 76608 142066 76664
rect 142122 76608 142127 76664
rect 141068 76606 142127 76608
rect 141068 76604 141074 76606
rect 142061 76603 142127 76606
rect 142337 76666 142403 76669
rect 142654 76666 142660 76668
rect 142337 76664 142660 76666
rect 142337 76608 142342 76664
rect 142398 76608 142660 76664
rect 142337 76606 142660 76608
rect 142337 76603 142403 76606
rect 142654 76604 142660 76606
rect 142724 76604 142730 76668
rect 143942 76604 143948 76668
rect 144012 76666 144018 76668
rect 144545 76666 144611 76669
rect 144012 76664 144611 76666
rect 144012 76608 144550 76664
rect 144606 76608 144611 76664
rect 144012 76606 144611 76608
rect 144012 76604 144018 76606
rect 144545 76603 144611 76606
rect 146518 76604 146524 76668
rect 146588 76666 146594 76668
rect 146661 76666 146727 76669
rect 146588 76664 146727 76666
rect 146588 76608 146666 76664
rect 146722 76608 146727 76664
rect 146588 76606 146727 76608
rect 146588 76604 146594 76606
rect 146661 76603 146727 76606
rect 148041 76666 148107 76669
rect 148174 76666 148180 76668
rect 148041 76664 148180 76666
rect 148041 76608 148046 76664
rect 148102 76608 148180 76664
rect 148041 76606 148180 76608
rect 148041 76603 148107 76606
rect 148174 76604 148180 76606
rect 148244 76604 148250 76668
rect 149646 76604 149652 76668
rect 149716 76666 149722 76668
rect 150065 76666 150131 76669
rect 149716 76664 150131 76666
rect 149716 76608 150070 76664
rect 150126 76608 150131 76664
rect 149716 76606 150131 76608
rect 149716 76604 149722 76606
rect 150065 76603 150131 76606
rect 181437 76666 181503 76669
rect 535453 76666 535519 76669
rect 181437 76664 535519 76666
rect 181437 76608 181442 76664
rect 181498 76608 535458 76664
rect 535514 76608 535519 76664
rect 181437 76606 535519 76608
rect 181437 76603 181503 76606
rect 535453 76603 535519 76606
rect 115933 76530 115999 76533
rect 139342 76530 139348 76532
rect 115933 76528 139348 76530
rect 115933 76472 115938 76528
rect 115994 76472 139348 76528
rect 115933 76470 139348 76472
rect 115933 76467 115999 76470
rect 139342 76468 139348 76470
rect 139412 76468 139418 76532
rect 174997 76530 175063 76533
rect 549253 76530 549319 76533
rect 174997 76528 549319 76530
rect 174997 76472 175002 76528
rect 175058 76472 549258 76528
rect 549314 76472 549319 76528
rect 174997 76470 549319 76472
rect 174997 76467 175063 76470
rect 549253 76467 549319 76470
rect 172237 76394 172303 76397
rect 181437 76394 181503 76397
rect 172237 76392 181503 76394
rect 172237 76336 172242 76392
rect 172298 76336 181442 76392
rect 181498 76336 181503 76392
rect 172237 76334 181503 76336
rect 172237 76331 172303 76334
rect 181437 76331 181503 76334
rect 156822 76196 156828 76260
rect 156892 76258 156898 76260
rect 158253 76258 158319 76261
rect 156892 76256 158319 76258
rect 156892 76200 158258 76256
rect 158314 76200 158319 76256
rect 156892 76198 158319 76200
rect 156892 76196 156898 76198
rect 158253 76195 158319 76198
rect 148777 76122 148843 76125
rect 149421 76124 149487 76125
rect 148910 76122 148916 76124
rect 148777 76120 148916 76122
rect 148777 76064 148782 76120
rect 148838 76064 148916 76120
rect 148777 76062 148916 76064
rect 148777 76059 148843 76062
rect 148910 76060 148916 76062
rect 148980 76060 148986 76124
rect 149421 76122 149468 76124
rect 149376 76120 149468 76122
rect 149376 76064 149426 76120
rect 149376 76062 149468 76064
rect 149421 76060 149468 76062
rect 149532 76060 149538 76124
rect 152774 76060 152780 76124
rect 152844 76122 152850 76124
rect 153101 76122 153167 76125
rect 152844 76120 153167 76122
rect 152844 76064 153106 76120
rect 153162 76064 153167 76120
rect 152844 76062 153167 76064
rect 152844 76060 152850 76062
rect 149421 76059 149487 76060
rect 153101 76059 153167 76062
rect 156638 76060 156644 76124
rect 156708 76122 156714 76124
rect 157149 76122 157215 76125
rect 156708 76120 157215 76122
rect 156708 76064 157154 76120
rect 157210 76064 157215 76120
rect 156708 76062 157215 76064
rect 156708 76060 156714 76062
rect 157149 76059 157215 76062
rect 171358 76060 171364 76124
rect 171428 76122 171434 76124
rect 177062 76122 177068 76124
rect 171428 76062 177068 76122
rect 171428 76060 171434 76062
rect 177062 76060 177068 76062
rect 177132 76060 177138 76124
rect 148542 75924 148548 75988
rect 148612 75986 148618 75988
rect 148869 75986 148935 75989
rect 148612 75984 148935 75986
rect 148612 75928 148874 75984
rect 148930 75928 148935 75984
rect 148612 75926 148935 75928
rect 148612 75924 148618 75926
rect 148869 75923 148935 75926
rect 149094 75924 149100 75988
rect 149164 75986 149170 75988
rect 149697 75986 149763 75989
rect 149164 75984 149763 75986
rect 149164 75928 149702 75984
rect 149758 75928 149763 75984
rect 149164 75926 149763 75928
rect 149164 75924 149170 75926
rect 149697 75923 149763 75926
rect 149973 75988 150039 75989
rect 149973 75984 150020 75988
rect 150084 75986 150090 75988
rect 150709 75986 150775 75989
rect 151118 75986 151124 75988
rect 149973 75928 149978 75984
rect 149973 75924 150020 75928
rect 150084 75926 150130 75986
rect 150709 75984 151124 75986
rect 150709 75928 150714 75984
rect 150770 75928 151124 75984
rect 150709 75926 151124 75928
rect 150084 75924 150090 75926
rect 149973 75923 150039 75924
rect 150709 75923 150775 75926
rect 151118 75924 151124 75926
rect 151188 75924 151194 75988
rect 151486 75924 151492 75988
rect 151556 75986 151562 75988
rect 151629 75986 151695 75989
rect 152181 75988 152247 75989
rect 152181 75986 152228 75988
rect 151556 75984 151695 75986
rect 151556 75928 151634 75984
rect 151690 75928 151695 75984
rect 151556 75926 151695 75928
rect 152136 75984 152228 75986
rect 152136 75928 152186 75984
rect 152136 75926 152228 75928
rect 151556 75924 151562 75926
rect 151629 75923 151695 75926
rect 152181 75924 152228 75926
rect 152292 75924 152298 75988
rect 152825 75986 152891 75989
rect 152958 75986 152964 75988
rect 152825 75984 152964 75986
rect 152825 75928 152830 75984
rect 152886 75928 152964 75984
rect 152825 75926 152964 75928
rect 152181 75923 152247 75924
rect 152825 75923 152891 75926
rect 152958 75924 152964 75926
rect 153028 75924 153034 75988
rect 153561 75986 153627 75989
rect 153694 75986 153700 75988
rect 153561 75984 153700 75986
rect 153561 75928 153566 75984
rect 153622 75928 153700 75984
rect 153561 75926 153700 75928
rect 153561 75923 153627 75926
rect 153694 75924 153700 75926
rect 153764 75924 153770 75988
rect 154246 75924 154252 75988
rect 154316 75986 154322 75988
rect 154481 75986 154547 75989
rect 154316 75984 154547 75986
rect 154316 75928 154486 75984
rect 154542 75928 154547 75984
rect 154316 75926 154547 75928
rect 154316 75924 154322 75926
rect 154481 75923 154547 75926
rect 154614 75924 154620 75988
rect 154684 75986 154690 75988
rect 156965 75986 157031 75989
rect 154684 75984 157031 75986
rect 154684 75928 156970 75984
rect 157026 75928 157031 75984
rect 154684 75926 157031 75928
rect 154684 75924 154690 75926
rect 156965 75923 157031 75926
rect 168649 75986 168715 75989
rect 169150 75986 169156 75988
rect 168649 75984 169156 75986
rect 168649 75928 168654 75984
rect 168710 75928 169156 75984
rect 168649 75926 169156 75928
rect 168649 75923 168715 75926
rect 169150 75924 169156 75926
rect 169220 75924 169226 75988
rect 170070 75924 170076 75988
rect 170140 75986 170146 75988
rect 170213 75986 170279 75989
rect 170857 75988 170923 75989
rect 170806 75986 170812 75988
rect 170140 75984 170279 75986
rect 170140 75928 170218 75984
rect 170274 75928 170279 75984
rect 170140 75926 170279 75928
rect 170766 75926 170812 75986
rect 170876 75984 170923 75988
rect 170918 75928 170923 75984
rect 170140 75924 170146 75926
rect 170213 75923 170279 75926
rect 170806 75924 170812 75926
rect 170876 75924 170923 75928
rect 171542 75924 171548 75988
rect 171612 75986 171618 75988
rect 171777 75986 171843 75989
rect 171612 75984 171843 75986
rect 171612 75928 171782 75984
rect 171838 75928 171843 75984
rect 171612 75926 171843 75928
rect 171612 75924 171618 75926
rect 170857 75923 170923 75924
rect 171777 75923 171843 75926
rect 175457 75986 175523 75989
rect 175958 75986 175964 75988
rect 175457 75984 175964 75986
rect 175457 75928 175462 75984
rect 175518 75928 175964 75984
rect 175457 75926 175964 75928
rect 175457 75923 175523 75926
rect 175958 75924 175964 75926
rect 176028 75924 176034 75988
rect 176610 75926 177130 75986
rect 132585 75850 132651 75853
rect 133270 75850 133276 75852
rect 132585 75848 133276 75850
rect 132585 75792 132590 75848
rect 132646 75792 133276 75848
rect 132585 75790 133276 75792
rect 132585 75787 132651 75790
rect 133270 75788 133276 75790
rect 133340 75788 133346 75852
rect 144678 75788 144684 75852
rect 144748 75850 144754 75852
rect 176610 75850 176670 75926
rect 144748 75790 176670 75850
rect 177070 75850 177130 75926
rect 177389 75850 177455 75853
rect 177070 75848 177455 75850
rect 177070 75792 177394 75848
rect 177450 75792 177455 75848
rect 177070 75790 177455 75792
rect 144748 75788 144754 75790
rect 177389 75787 177455 75790
rect 155677 75714 155743 75717
rect 272885 75714 272951 75717
rect 155677 75712 272951 75714
rect 155677 75656 155682 75712
rect 155738 75656 272890 75712
rect 272946 75656 272951 75712
rect 155677 75654 272951 75656
rect 155677 75651 155743 75654
rect 272885 75651 272951 75654
rect 156781 75578 156847 75581
rect 305637 75578 305703 75581
rect 156781 75576 305703 75578
rect 156781 75520 156786 75576
rect 156842 75520 305642 75576
rect 305698 75520 305703 75576
rect 156781 75518 305703 75520
rect 156781 75515 156847 75518
rect 305637 75515 305703 75518
rect 80053 75442 80119 75445
rect 136582 75442 136588 75444
rect 80053 75440 136588 75442
rect 80053 75384 80058 75440
rect 80114 75384 136588 75440
rect 80053 75382 136588 75384
rect 80053 75379 80119 75382
rect 136582 75380 136588 75382
rect 136652 75380 136658 75444
rect 156873 75442 156939 75445
rect 310237 75442 310303 75445
rect 156873 75440 310303 75442
rect 156873 75384 156878 75440
rect 156934 75384 310242 75440
rect 310298 75384 310303 75440
rect 156873 75382 310303 75384
rect 156873 75379 156939 75382
rect 310237 75379 310303 75382
rect 46933 75306 46999 75309
rect 132401 75306 132467 75309
rect 46933 75304 132467 75306
rect 46933 75248 46938 75304
rect 46994 75248 132406 75304
rect 132462 75248 132467 75304
rect 46933 75246 132467 75248
rect 46933 75243 46999 75246
rect 132401 75243 132467 75246
rect 175089 75304 175155 75309
rect 175089 75248 175094 75304
rect 175150 75248 175155 75304
rect 175089 75243 175155 75248
rect 175365 75306 175431 75309
rect 547873 75306 547939 75309
rect 175365 75304 547939 75306
rect 175365 75248 175370 75304
rect 175426 75248 547878 75304
rect 547934 75248 547939 75304
rect 175365 75246 547939 75248
rect 175365 75243 175431 75246
rect 547873 75243 547939 75246
rect 6913 75170 6979 75173
rect 126881 75170 126947 75173
rect 6913 75168 126947 75170
rect 6913 75112 6918 75168
rect 6974 75112 126886 75168
rect 126942 75112 126947 75168
rect 6913 75110 126947 75112
rect 175092 75170 175152 75243
rect 571333 75170 571399 75173
rect 175092 75168 571399 75170
rect 175092 75112 571338 75168
rect 571394 75112 571399 75168
rect 175092 75110 571399 75112
rect 6913 75107 6979 75110
rect 126881 75107 126947 75110
rect 571333 75107 571399 75110
rect 155902 74972 155908 75036
rect 155972 75034 155978 75036
rect 179413 75034 179479 75037
rect 155972 75032 179479 75034
rect 155972 74976 179418 75032
rect 179474 74976 179479 75032
rect 155972 74974 179479 74976
rect 155972 74972 155978 74974
rect 179413 74971 179479 74974
rect 160001 74898 160067 74901
rect 178953 74898 179019 74901
rect 160001 74896 179019 74898
rect 160001 74840 160006 74896
rect 160062 74840 178958 74896
rect 179014 74840 179019 74896
rect 160001 74838 179019 74840
rect 160001 74835 160067 74838
rect 178953 74835 179019 74838
rect 160870 74564 160876 74628
rect 160940 74626 160946 74628
rect 161422 74626 161428 74628
rect 160940 74566 161428 74626
rect 160940 74564 160946 74566
rect 161422 74564 161428 74566
rect 161492 74564 161498 74628
rect 157006 74292 157012 74356
rect 157076 74354 157082 74356
rect 157609 74354 157675 74357
rect 157076 74352 157675 74354
rect 157076 74296 157614 74352
rect 157670 74296 157675 74352
rect 157076 74294 157675 74296
rect 157076 74292 157082 74294
rect 157609 74291 157675 74294
rect 161238 74156 161244 74220
rect 161308 74218 161314 74220
rect 178861 74218 178927 74221
rect 161308 74216 178927 74218
rect 161308 74160 178866 74216
rect 178922 74160 178927 74216
rect 161308 74158 178927 74160
rect 161308 74156 161314 74158
rect 178861 74155 178927 74158
rect 150249 74082 150315 74085
rect 251173 74082 251239 74085
rect 150249 74080 251239 74082
rect 150249 74024 150254 74080
rect 150310 74024 251178 74080
rect 251234 74024 251239 74080
rect 150249 74022 251239 74024
rect 150249 74019 150315 74022
rect 251173 74019 251239 74022
rect 157241 73946 157307 73949
rect 295333 73946 295399 73949
rect 157241 73944 295399 73946
rect 157241 73888 157246 73944
rect 157302 73888 295338 73944
rect 295394 73888 295399 73944
rect 157241 73886 295399 73888
rect 157241 73883 157307 73886
rect 295333 73883 295399 73886
rect 64873 73810 64939 73813
rect 135846 73810 135852 73812
rect 64873 73808 135852 73810
rect 64873 73752 64878 73808
rect 64934 73752 135852 73808
rect 64873 73750 135852 73752
rect 64873 73747 64939 73750
rect 135846 73748 135852 73750
rect 135916 73748 135922 73812
rect 156454 73748 156460 73812
rect 156524 73810 156530 73812
rect 157609 73810 157675 73813
rect 156524 73808 157675 73810
rect 156524 73752 157614 73808
rect 157670 73752 157675 73808
rect 156524 73750 157675 73752
rect 156524 73748 156530 73750
rect 157609 73747 157675 73750
rect 158621 73810 158687 73813
rect 318149 73810 318215 73813
rect 158621 73808 318215 73810
rect 158621 73752 158626 73808
rect 158682 73752 318154 73808
rect 318210 73752 318215 73808
rect 158621 73750 318215 73752
rect 158621 73747 158687 73750
rect 318149 73747 318215 73750
rect 174486 73476 174492 73540
rect 174556 73538 174562 73540
rect 176469 73538 176535 73541
rect 174556 73536 176535 73538
rect 174556 73480 176474 73536
rect 176530 73480 176535 73536
rect 174556 73478 176535 73480
rect 174556 73476 174562 73478
rect 176469 73475 176535 73478
rect 131113 73268 131179 73269
rect 131062 73204 131068 73268
rect 131132 73266 131179 73268
rect 131132 73264 131224 73266
rect 131174 73208 131224 73264
rect 131132 73206 131224 73208
rect 131132 73204 131179 73206
rect 131113 73203 131179 73204
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 97993 72722 98059 72725
rect 138422 72722 138428 72724
rect 97993 72720 138428 72722
rect 97993 72664 97998 72720
rect 98054 72664 138428 72720
rect 97993 72662 138428 72664
rect 97993 72659 98059 72662
rect 138422 72660 138428 72662
rect 138492 72660 138498 72724
rect 27613 72586 27679 72589
rect 130745 72586 130811 72589
rect 27613 72584 130811 72586
rect 27613 72528 27618 72584
rect 27674 72528 130750 72584
rect 130806 72528 130811 72584
rect 27613 72526 130811 72528
rect 27613 72523 27679 72526
rect 130745 72523 130811 72526
rect 158294 72524 158300 72588
rect 158364 72586 158370 72588
rect 289169 72586 289235 72589
rect 158364 72584 289235 72586
rect 158364 72528 289174 72584
rect 289230 72528 289235 72584
rect 158364 72526 289235 72528
rect 158364 72524 158370 72526
rect 289169 72523 289235 72526
rect 8293 72450 8359 72453
rect 131614 72450 131620 72452
rect 8293 72448 131620 72450
rect 8293 72392 8298 72448
rect 8354 72392 131620 72448
rect 8293 72390 131620 72392
rect 8293 72387 8359 72390
rect 131614 72388 131620 72390
rect 131684 72388 131690 72452
rect 168046 72388 168052 72452
rect 168116 72450 168122 72452
rect 445477 72450 445543 72453
rect 168116 72448 445543 72450
rect 168116 72392 445482 72448
rect 445538 72392 445543 72448
rect 168116 72390 445543 72392
rect 168116 72388 168122 72390
rect 445477 72387 445543 72390
rect -960 71634 480 71724
rect 158110 71708 158116 71772
rect 158180 71770 158186 71772
rect 261569 71770 261635 71773
rect 158180 71768 261635 71770
rect 158180 71712 261574 71768
rect 261630 71712 261635 71768
rect 158180 71710 261635 71712
rect 158180 71708 158186 71710
rect 261569 71707 261635 71710
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 156638 71572 156644 71636
rect 156708 71634 156714 71636
rect 280889 71634 280955 71637
rect 156708 71632 280955 71634
rect 156708 71576 280894 71632
rect 280950 71576 280955 71632
rect 156708 71574 280955 71576
rect 156708 71572 156714 71574
rect 280889 71571 280955 71574
rect 158846 71436 158852 71500
rect 158916 71498 158922 71500
rect 310421 71498 310487 71501
rect 158916 71496 310487 71498
rect 158916 71440 310426 71496
rect 310482 71440 310487 71496
rect 158916 71438 310487 71440
rect 158916 71436 158922 71438
rect 310421 71435 310487 71438
rect 161422 71300 161428 71364
rect 161492 71362 161498 71364
rect 396073 71362 396139 71365
rect 161492 71360 396139 71362
rect 161492 71304 396078 71360
rect 396134 71304 396139 71360
rect 161492 71302 396139 71304
rect 161492 71300 161498 71302
rect 396073 71299 396139 71302
rect 169702 71164 169708 71228
rect 169772 71226 169778 71228
rect 500953 71226 501019 71229
rect 169772 71224 501019 71226
rect 169772 71168 500958 71224
rect 501014 71168 501019 71224
rect 169772 71166 501019 71168
rect 169772 71164 169778 71166
rect 500953 71163 501019 71166
rect 170622 71028 170628 71092
rect 170692 71090 170698 71092
rect 518893 71090 518959 71093
rect 170692 71088 518959 71090
rect 170692 71032 518898 71088
rect 518954 71032 518959 71088
rect 170692 71030 518959 71032
rect 170692 71028 170698 71030
rect 518893 71027 518959 71030
rect 167678 69532 167684 69596
rect 167748 69594 167754 69596
rect 475377 69594 475443 69597
rect 167748 69592 475443 69594
rect 167748 69536 475382 69592
rect 475438 69536 475443 69592
rect 167748 69534 475443 69536
rect 167748 69532 167754 69534
rect 475377 69531 475443 69534
rect 144310 68444 144316 68508
rect 144380 68506 144386 68508
rect 179413 68506 179479 68509
rect 144380 68504 179479 68506
rect 144380 68448 179418 68504
rect 179474 68448 179479 68504
rect 144380 68446 179479 68448
rect 144380 68444 144386 68446
rect 179413 68443 179479 68446
rect 158478 68308 158484 68372
rect 158548 68370 158554 68372
rect 303245 68370 303311 68373
rect 158548 68368 303311 68370
rect 158548 68312 303250 68368
rect 303306 68312 303311 68368
rect 158548 68310 303311 68312
rect 158548 68308 158554 68310
rect 303245 68307 303311 68310
rect 167862 68172 167868 68236
rect 167932 68234 167938 68236
rect 439497 68234 439563 68237
rect 167932 68232 439563 68234
rect 167932 68176 439502 68232
rect 439558 68176 439563 68232
rect 167932 68174 439563 68176
rect 167932 68172 167938 68174
rect 439497 68171 439563 68174
rect 144494 66812 144500 66876
rect 144564 66874 144570 66876
rect 182173 66874 182239 66877
rect 144564 66872 182239 66874
rect 144564 66816 182178 66872
rect 182234 66816 182239 66872
rect 144564 66814 182239 66816
rect 144564 66812 144570 66814
rect 182173 66811 182239 66814
rect 145230 63004 145236 63068
rect 145300 63066 145306 63068
rect 200113 63066 200179 63069
rect 145300 63064 200179 63066
rect 145300 63008 200118 63064
rect 200174 63008 200179 63064
rect 145300 63006 200179 63008
rect 145300 63004 145306 63006
rect 200113 63003 200179 63006
rect 174854 62868 174860 62932
rect 174924 62930 174930 62932
rect 572713 62930 572779 62933
rect 174924 62928 572779 62930
rect 174924 62872 572718 62928
rect 572774 62872 572779 62928
rect 174924 62870 572779 62872
rect 174924 62868 174930 62870
rect 572713 62867 572779 62870
rect 176142 62732 176148 62796
rect 176212 62794 176218 62796
rect 581085 62794 581151 62797
rect 176212 62792 581151 62794
rect 176212 62736 581090 62792
rect 581146 62736 581151 62792
rect 176212 62734 581151 62736
rect 176212 62732 176218 62734
rect 581085 62731 581151 62734
rect 171910 61508 171916 61572
rect 171980 61570 171986 61572
rect 536833 61570 536899 61573
rect 171980 61568 536899 61570
rect 171980 61512 536838 61568
rect 536894 61512 536899 61568
rect 171980 61510 536899 61512
rect 171980 61508 171986 61510
rect 536833 61507 536899 61510
rect 176326 61372 176332 61436
rect 176396 61434 176402 61436
rect 575473 61434 575539 61437
rect 176396 61432 575539 61434
rect 176396 61376 575478 61432
rect 575534 61376 575539 61432
rect 176396 61374 575539 61376
rect 176396 61372 176402 61374
rect 575473 61371 575539 61374
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 144126 57156 144132 57220
rect 144196 57218 144202 57220
rect 183553 57218 183619 57221
rect 144196 57216 183619 57218
rect 144196 57160 183558 57216
rect 183614 57160 183619 57216
rect 144196 57158 183619 57160
rect 144196 57156 144202 57158
rect 183553 57155 183619 57158
rect 161054 48860 161060 48924
rect 161124 48922 161130 48924
rect 394693 48922 394759 48925
rect 161124 48920 394759 48922
rect 161124 48864 394698 48920
rect 394754 48864 394759 48920
rect 161124 48862 394759 48864
rect 161124 48860 161130 48862
rect 394693 48859 394759 48862
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 176510 46140 176516 46204
rect 176580 46202 176586 46204
rect 576853 46202 576919 46205
rect 176580 46200 576919 46202
rect 176580 46144 576858 46200
rect 576914 46144 576919 46200
rect 583520 46188 584960 46278
rect 176580 46142 576919 46144
rect 176580 46140 176586 46142
rect 576853 46139 576919 46142
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 11145 35186 11211 35189
rect 131246 35186 131252 35188
rect 11145 35184 131252 35186
rect 11145 35128 11150 35184
rect 11206 35128 131252 35184
rect 11145 35126 131252 35128
rect 11145 35123 11211 35126
rect 131246 35124 131252 35126
rect 131316 35124 131322 35188
rect 147070 34172 147076 34236
rect 147140 34234 147146 34236
rect 216673 34234 216739 34237
rect 147140 34232 216739 34234
rect 147140 34176 216678 34232
rect 216734 34176 216739 34232
rect 147140 34174 216739 34176
rect 147140 34172 147146 34174
rect 216673 34171 216739 34174
rect 163446 34036 163452 34100
rect 163516 34098 163522 34100
rect 429193 34098 429259 34101
rect 163516 34096 429259 34098
rect 163516 34040 429198 34096
rect 429254 34040 429259 34096
rect 163516 34038 429259 34040
rect 163516 34036 163522 34038
rect 429193 34035 429259 34038
rect 163262 33900 163268 33964
rect 163332 33962 163338 33964
rect 432045 33962 432111 33965
rect 163332 33960 432111 33962
rect 163332 33904 432050 33960
rect 432106 33904 432111 33960
rect 163332 33902 432111 33904
rect 163332 33900 163338 33902
rect 432045 33899 432111 33902
rect 173566 33764 173572 33828
rect 173636 33826 173642 33828
rect 556153 33826 556219 33829
rect 173636 33824 556219 33826
rect 173636 33768 556158 33824
rect 556214 33768 556219 33824
rect 173636 33766 556219 33768
rect 173636 33764 173642 33766
rect 556153 33763 556219 33766
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 163630 31316 163636 31380
rect 163700 31378 163706 31380
rect 430573 31378 430639 31381
rect 163700 31376 430639 31378
rect 163700 31320 430578 31376
rect 430634 31320 430639 31376
rect 163700 31318 430639 31320
rect 163700 31316 163706 31318
rect 430573 31315 430639 31318
rect 166206 31180 166212 31244
rect 166276 31242 166282 31244
rect 465073 31242 465139 31245
rect 166276 31240 465139 31242
rect 166276 31184 465078 31240
rect 465134 31184 465139 31240
rect 166276 31182 465139 31184
rect 166276 31180 166282 31182
rect 465073 31179 465139 31182
rect 167494 31044 167500 31108
rect 167564 31106 167570 31108
rect 483013 31106 483079 31109
rect 167564 31104 483079 31106
rect 167564 31048 483018 31104
rect 483074 31048 483079 31104
rect 167564 31046 483079 31048
rect 167564 31044 167570 31046
rect 483013 31043 483079 31046
rect 173750 30908 173756 30972
rect 173820 30970 173826 30972
rect 554773 30970 554839 30973
rect 173820 30968 554839 30970
rect 173820 30912 554778 30968
rect 554834 30912 554839 30968
rect 173820 30910 554839 30912
rect 173820 30908 173826 30910
rect 554773 30907 554839 30910
rect 151302 28460 151308 28524
rect 151372 28522 151378 28524
rect 292573 28522 292639 28525
rect 151372 28520 292639 28522
rect 151372 28464 292578 28520
rect 292634 28464 292639 28520
rect 151372 28462 292639 28464
rect 151372 28460 151378 28462
rect 292573 28459 292639 28462
rect 166390 28324 166396 28388
rect 166460 28386 166466 28388
rect 466453 28386 466519 28389
rect 166460 28384 466519 28386
rect 166460 28328 466458 28384
rect 466514 28328 466519 28384
rect 166460 28326 466519 28328
rect 166460 28324 166466 28326
rect 466453 28323 466519 28326
rect 171777 28250 171843 28253
rect 531313 28250 531379 28253
rect 171777 28248 531379 28250
rect 171777 28192 171782 28248
rect 171838 28192 531318 28248
rect 531374 28192 531379 28248
rect 171777 28190 531379 28192
rect 171777 28187 171843 28190
rect 531313 28187 531379 28190
rect 145414 25468 145420 25532
rect 145484 25530 145490 25532
rect 201585 25530 201651 25533
rect 145484 25528 201651 25530
rect 145484 25472 201590 25528
rect 201646 25472 201651 25528
rect 145484 25470 201651 25472
rect 145484 25468 145490 25470
rect 201585 25467 201651 25470
rect 170806 24244 170812 24308
rect 170876 24306 170882 24308
rect 517513 24306 517579 24309
rect 170876 24304 517579 24306
rect 170876 24248 517518 24304
rect 517574 24248 517579 24304
rect 170876 24246 517579 24248
rect 170876 24244 170882 24246
rect 517513 24243 517579 24246
rect 174670 24108 174676 24172
rect 174740 24170 174746 24172
rect 569953 24170 570019 24173
rect 174740 24168 570019 24170
rect 174740 24112 569958 24168
rect 570014 24112 570019 24168
rect 174740 24110 570019 24112
rect 174740 24108 174746 24110
rect 569953 24107 570019 24110
rect 147254 23292 147260 23356
rect 147324 23354 147330 23356
rect 215293 23354 215359 23357
rect 147324 23352 215359 23354
rect 147324 23296 215298 23352
rect 215354 23296 215359 23352
rect 147324 23294 215359 23296
rect 147324 23292 147330 23294
rect 215293 23291 215359 23294
rect 152406 23156 152412 23220
rect 152476 23218 152482 23220
rect 284293 23218 284359 23221
rect 152476 23216 284359 23218
rect 152476 23160 284298 23216
rect 284354 23160 284359 23216
rect 152476 23158 284359 23160
rect 152476 23156 152482 23158
rect 284293 23155 284359 23158
rect 140630 23020 140636 23084
rect 140700 23082 140706 23084
rect 287053 23082 287119 23085
rect 140700 23080 287119 23082
rect 140700 23024 287058 23080
rect 287114 23024 287119 23080
rect 140700 23022 287119 23024
rect 140700 23020 140706 23022
rect 287053 23019 287119 23022
rect 170254 22884 170260 22948
rect 170324 22946 170330 22948
rect 516133 22946 516199 22949
rect 170324 22944 516199 22946
rect 170324 22888 516138 22944
rect 516194 22888 516199 22944
rect 170324 22886 516199 22888
rect 170324 22884 170330 22886
rect 516133 22883 516199 22886
rect 170990 22748 170996 22812
rect 171060 22810 171066 22812
rect 520273 22810 520339 22813
rect 171060 22808 520339 22810
rect 171060 22752 520278 22808
rect 520334 22752 520339 22808
rect 171060 22750 520339 22752
rect 171060 22748 171066 22750
rect 520273 22747 520339 22750
rect 60733 22674 60799 22677
rect 135662 22674 135668 22676
rect 60733 22672 135668 22674
rect 60733 22616 60738 22672
rect 60794 22616 135668 22672
rect 60733 22614 135668 22616
rect 60733 22611 60799 22614
rect 135662 22612 135668 22614
rect 135732 22612 135738 22676
rect 172094 22612 172100 22676
rect 172164 22674 172170 22676
rect 538213 22674 538279 22677
rect 172164 22672 538279 22674
rect 172164 22616 538218 22672
rect 538274 22616 538279 22672
rect 172164 22614 538279 22616
rect 172164 22612 172170 22614
rect 538213 22611 538279 22614
rect 169518 21252 169524 21316
rect 169588 21314 169594 21316
rect 502333 21314 502399 21317
rect 169588 21312 502399 21314
rect 169588 21256 502338 21312
rect 502394 21256 502399 21312
rect 169588 21254 502399 21256
rect 169588 21252 169594 21254
rect 502333 21251 502399 21254
rect 145598 20436 145604 20500
rect 145668 20498 145674 20500
rect 241513 20498 241579 20501
rect 145668 20496 241579 20498
rect 145668 20440 241518 20496
rect 241574 20440 241579 20496
rect 145668 20438 241579 20440
rect 145668 20436 145674 20438
rect 241513 20435 241579 20438
rect 139158 20300 139164 20364
rect 139228 20362 139234 20364
rect 266353 20362 266419 20365
rect 139228 20360 266419 20362
rect 139228 20304 266358 20360
rect 266414 20304 266419 20360
rect 139228 20302 266419 20304
rect 139228 20300 139234 20302
rect 266353 20299 266419 20302
rect 162342 20164 162348 20228
rect 162412 20226 162418 20228
rect 409873 20226 409939 20229
rect 162412 20224 409939 20226
rect 162412 20168 409878 20224
rect 409934 20168 409939 20224
rect 162412 20166 409939 20168
rect 162412 20164 162418 20166
rect 409873 20163 409939 20166
rect 162158 20028 162164 20092
rect 162228 20090 162234 20092
rect 414013 20090 414079 20093
rect 162228 20088 414079 20090
rect 162228 20032 414018 20088
rect 414074 20032 414079 20088
rect 162228 20030 414079 20032
rect 162228 20028 162234 20030
rect 414013 20027 414079 20030
rect 171726 19892 171732 19956
rect 171796 19954 171802 19956
rect 534073 19954 534139 19957
rect 171796 19952 534139 19954
rect 171796 19896 534078 19952
rect 534134 19896 534139 19952
rect 171796 19894 534139 19896
rect 171796 19892 171802 19894
rect 534073 19891 534139 19894
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 2957 19410 3023 19413
rect -960 19408 3023 19410
rect -960 19352 2962 19408
rect 3018 19352 3023 19408
rect -960 19350 3023 19352
rect -960 19260 480 19350
rect 2957 19347 3023 19350
rect 142838 18668 142844 18732
rect 142908 18730 142914 18732
rect 162945 18730 163011 18733
rect 142908 18728 163011 18730
rect 142908 18672 162950 18728
rect 163006 18672 163011 18728
rect 142908 18670 163011 18672
rect 142908 18668 142914 18670
rect 162945 18667 163011 18670
rect 148358 18532 148364 18596
rect 148428 18594 148434 18596
rect 234613 18594 234679 18597
rect 148428 18592 234679 18594
rect 148428 18536 234618 18592
rect 234674 18536 234679 18592
rect 148428 18534 234679 18536
rect 148428 18532 148434 18534
rect 234613 18531 234679 18534
rect 165286 17716 165292 17780
rect 165356 17778 165362 17780
rect 444373 17778 444439 17781
rect 165356 17776 444439 17778
rect 165356 17720 444378 17776
rect 444434 17720 444439 17776
rect 165356 17718 444439 17720
rect 165356 17716 165362 17718
rect 444373 17715 444439 17718
rect 165102 17580 165108 17644
rect 165172 17642 165178 17644
rect 445753 17642 445819 17645
rect 165172 17640 445819 17642
rect 165172 17584 445758 17640
rect 445814 17584 445819 17640
rect 165172 17582 445819 17584
rect 165172 17580 165178 17582
rect 445753 17579 445819 17582
rect 164918 17444 164924 17508
rect 164988 17506 164994 17508
rect 448513 17506 448579 17509
rect 164988 17504 448579 17506
rect 164988 17448 448518 17504
rect 448574 17448 448579 17504
rect 164988 17446 448579 17448
rect 164988 17444 164994 17446
rect 448513 17443 448579 17446
rect 166758 17308 166764 17372
rect 166828 17370 166834 17372
rect 463693 17370 463759 17373
rect 166828 17368 463759 17370
rect 166828 17312 463698 17368
rect 463754 17312 463759 17368
rect 166828 17310 463759 17312
rect 166828 17308 166834 17310
rect 463693 17307 463759 17310
rect 166574 17172 166580 17236
rect 166644 17234 166650 17236
rect 465165 17234 465231 17237
rect 166644 17232 465231 17234
rect 166644 17176 465170 17232
rect 465226 17176 465231 17232
rect 166644 17174 465231 17176
rect 166644 17172 166650 17174
rect 465165 17171 465231 17174
rect 152590 14452 152596 14516
rect 152660 14514 152666 14516
rect 286593 14514 286659 14517
rect 152660 14512 286659 14514
rect 152660 14456 286598 14512
rect 286654 14456 286659 14512
rect 152660 14454 286659 14456
rect 152660 14452 152666 14454
rect 286593 14451 286659 14454
rect 149646 12004 149652 12068
rect 149716 12066 149722 12068
rect 251265 12066 251331 12069
rect 149716 12064 251331 12066
rect 149716 12008 251270 12064
rect 251326 12008 251331 12064
rect 149716 12006 251331 12008
rect 149716 12004 149722 12006
rect 251265 12003 251331 12006
rect 151486 11868 151492 11932
rect 151556 11930 151562 11932
rect 272425 11930 272491 11933
rect 151556 11928 272491 11930
rect 151556 11872 272430 11928
rect 272486 11872 272491 11928
rect 151556 11870 272491 11872
rect 151556 11868 151562 11870
rect 272425 11867 272491 11870
rect 162526 11732 162532 11796
rect 162596 11794 162602 11796
rect 409137 11794 409203 11797
rect 162596 11792 409203 11794
rect 162596 11736 409142 11792
rect 409198 11736 409203 11792
rect 162596 11734 409203 11736
rect 162596 11732 162602 11734
rect 409137 11731 409203 11734
rect 114001 11658 114067 11661
rect 139526 11658 139532 11660
rect 114001 11656 139532 11658
rect 114001 11600 114006 11656
rect 114062 11600 139532 11656
rect 114001 11598 139532 11600
rect 114001 11595 114067 11598
rect 139526 11596 139532 11598
rect 139596 11596 139602 11660
rect 162710 11596 162716 11660
rect 162780 11658 162786 11660
rect 412633 11658 412699 11661
rect 162780 11656 412699 11658
rect 162780 11600 412638 11656
rect 412694 11600 412699 11656
rect 162780 11598 412699 11600
rect 162780 11596 162786 11598
rect 412633 11595 412699 11598
rect 95785 10434 95851 10437
rect 138238 10434 138244 10436
rect 95785 10432 138244 10434
rect 95785 10376 95790 10432
rect 95846 10376 138244 10432
rect 95785 10374 138244 10376
rect 95785 10371 95851 10374
rect 138238 10372 138244 10374
rect 138308 10372 138314 10436
rect 148542 10372 148548 10436
rect 148612 10434 148618 10436
rect 236545 10434 236611 10437
rect 148612 10432 236611 10434
rect 148612 10376 236550 10432
rect 236606 10376 236611 10432
rect 148612 10374 236611 10376
rect 148612 10372 148618 10374
rect 236545 10371 236611 10374
rect 78121 10298 78187 10301
rect 137502 10298 137508 10300
rect 78121 10296 137508 10298
rect 78121 10240 78126 10296
rect 78182 10240 137508 10296
rect 78121 10238 137508 10240
rect 78121 10235 78187 10238
rect 137502 10236 137508 10238
rect 137572 10236 137578 10300
rect 160686 10236 160692 10300
rect 160756 10298 160762 10300
rect 392577 10298 392643 10301
rect 160756 10296 392643 10298
rect 160756 10240 392582 10296
rect 392638 10240 392643 10296
rect 160756 10238 392643 10240
rect 160756 10236 160762 10238
rect 392577 10235 392643 10238
rect 153878 9148 153884 9212
rect 153948 9210 153954 9212
rect 303153 9210 303219 9213
rect 153948 9208 303219 9210
rect 153948 9152 303158 9208
rect 303214 9152 303219 9208
rect 153948 9150 303219 9152
rect 153948 9148 153954 9150
rect 303153 9147 303219 9150
rect 119889 9074 119955 9077
rect 139710 9074 139716 9076
rect 119889 9072 139716 9074
rect 119889 9016 119894 9072
rect 119950 9016 139716 9072
rect 119889 9014 139716 9016
rect 119889 9011 119955 9014
rect 139710 9012 139716 9014
rect 139780 9012 139786 9076
rect 154062 9012 154068 9076
rect 154132 9074 154138 9076
rect 306741 9074 306807 9077
rect 154132 9072 306807 9074
rect 154132 9016 306746 9072
rect 306802 9016 306807 9072
rect 154132 9014 306807 9016
rect 154132 9012 154138 9014
rect 306741 9011 306807 9014
rect 45461 8938 45527 8941
rect 134190 8938 134196 8940
rect 45461 8936 134196 8938
rect 45461 8880 45466 8936
rect 45522 8880 134196 8936
rect 45461 8878 134196 8880
rect 45461 8875 45527 8878
rect 134190 8876 134196 8878
rect 134260 8876 134266 8940
rect 154246 8876 154252 8940
rect 154316 8938 154322 8940
rect 307937 8938 308003 8941
rect 154316 8936 308003 8938
rect 154316 8880 307942 8936
rect 307998 8880 308003 8936
rect 154316 8878 308003 8880
rect 154316 8876 154322 8878
rect 307937 8875 308003 8878
rect 64321 7986 64387 7989
rect 135478 7986 135484 7988
rect 64321 7984 135484 7986
rect 64321 7928 64326 7984
rect 64382 7928 135484 7984
rect 64321 7926 135484 7928
rect 64321 7923 64387 7926
rect 135478 7924 135484 7926
rect 135548 7924 135554 7988
rect 63217 7850 63283 7853
rect 135294 7850 135300 7852
rect 63217 7848 135300 7850
rect 63217 7792 63222 7848
rect 63278 7792 135300 7848
rect 63217 7790 135300 7792
rect 63217 7787 63283 7790
rect 135294 7788 135300 7790
rect 135364 7788 135370 7852
rect 48957 7714 49023 7717
rect 134006 7714 134012 7716
rect 48957 7712 134012 7714
rect 48957 7656 48962 7712
rect 49018 7656 134012 7712
rect 48957 7654 134012 7656
rect 48957 7651 49023 7654
rect 134006 7652 134012 7654
rect 134076 7652 134082 7716
rect 44265 7578 44331 7581
rect 134374 7578 134380 7580
rect 44265 7576 134380 7578
rect 44265 7520 44270 7576
rect 44326 7520 134380 7576
rect 44265 7518 134380 7520
rect 44265 7515 44331 7518
rect 134374 7516 134380 7518
rect 134444 7516 134450 7580
rect 150014 6836 150020 6900
rect 150084 6898 150090 6900
rect 249977 6898 250043 6901
rect 150084 6896 250043 6898
rect 150084 6840 249982 6896
rect 250038 6840 250043 6896
rect 150084 6838 250043 6840
rect 150084 6836 150090 6838
rect 249977 6835 250043 6838
rect 149830 6700 149836 6764
rect 149900 6762 149906 6764
rect 253473 6762 253539 6765
rect 149900 6760 253539 6762
rect 149900 6704 253478 6760
rect 253534 6704 253539 6760
rect 149900 6702 253539 6704
rect 149900 6700 149906 6702
rect 253473 6699 253539 6702
rect -960 6490 480 6580
rect 151670 6564 151676 6628
rect 151740 6626 151746 6628
rect 271229 6626 271295 6629
rect 151740 6624 271295 6626
rect 151740 6568 271234 6624
rect 271290 6568 271295 6624
rect 151740 6566 271295 6568
rect 151740 6564 151746 6566
rect 271229 6563 271295 6566
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 88885 6490 88951 6493
rect 131062 6490 131068 6492
rect 88885 6488 131068 6490
rect 88885 6432 88890 6488
rect 88946 6432 131068 6488
rect 88885 6430 131068 6432
rect 88885 6427 88951 6430
rect 131062 6428 131068 6430
rect 131132 6428 131138 6492
rect 152958 6428 152964 6492
rect 153028 6490 153034 6492
rect 285397 6490 285463 6493
rect 153028 6488 285463 6490
rect 153028 6432 285402 6488
rect 285458 6432 285463 6488
rect 583520 6476 584960 6566
rect 153028 6430 285463 6432
rect 153028 6428 153034 6430
rect 285397 6427 285463 6430
rect 26509 6354 26575 6357
rect 133086 6354 133092 6356
rect 26509 6352 133092 6354
rect 26509 6296 26514 6352
rect 26570 6296 133092 6352
rect 26509 6294 133092 6296
rect 26509 6291 26575 6294
rect 133086 6292 133092 6294
rect 133156 6292 133162 6356
rect 152774 6292 152780 6356
rect 152844 6354 152850 6356
rect 288985 6354 289051 6357
rect 152844 6352 289051 6354
rect 152844 6296 288990 6352
rect 289046 6296 289051 6352
rect 152844 6294 289051 6296
rect 152844 6292 152850 6294
rect 288985 6291 289051 6294
rect 25313 6218 25379 6221
rect 133270 6218 133276 6220
rect 25313 6216 133276 6218
rect 25313 6160 25318 6216
rect 25374 6160 133276 6216
rect 25313 6158 133276 6160
rect 25313 6155 25379 6158
rect 133270 6156 133276 6158
rect 133340 6156 133346 6220
rect 165470 6156 165476 6220
rect 165540 6218 165546 6220
rect 449801 6218 449867 6221
rect 165540 6216 449867 6218
rect 165540 6160 449806 6216
rect 449862 6160 449867 6216
rect 165540 6158 449867 6160
rect 165540 6156 165546 6158
rect 449801 6155 449867 6158
rect 147438 6020 147444 6084
rect 147508 6082 147514 6084
rect 218145 6082 218211 6085
rect 147508 6080 218211 6082
rect 147508 6024 218150 6080
rect 218206 6024 218211 6080
rect 147508 6022 218211 6024
rect 147508 6020 147514 6022
rect 218145 6019 218211 6022
rect 143022 4932 143028 4996
rect 143092 4994 143098 4996
rect 162485 4994 162551 4997
rect 143092 4992 162551 4994
rect 143092 4936 162490 4992
rect 162546 4936 162551 4992
rect 143092 4934 162551 4936
rect 143092 4932 143098 4934
rect 162485 4931 162551 4934
rect 143206 4796 143212 4860
rect 143276 4858 143282 4860
rect 166073 4858 166139 4861
rect 143276 4856 166139 4858
rect 143276 4800 166078 4856
rect 166134 4800 166139 4856
rect 143276 4798 166139 4800
rect 143276 4796 143282 4798
rect 166073 4795 166139 4798
rect 148726 3980 148732 4044
rect 148796 4042 148802 4044
rect 232221 4042 232287 4045
rect 148796 4040 232287 4042
rect 148796 3984 232226 4040
rect 232282 3984 232287 4040
rect 148796 3982 232287 3984
rect 148796 3980 148802 3982
rect 232221 3979 232287 3982
rect 148910 3844 148916 3908
rect 148980 3906 148986 3908
rect 235809 3906 235875 3909
rect 148980 3904 235875 3906
rect 148980 3848 235814 3904
rect 235870 3848 235875 3904
rect 148980 3846 235875 3848
rect 148980 3844 148986 3846
rect 235809 3843 235875 3846
rect 150065 3770 150131 3773
rect 242985 3770 243051 3773
rect 150065 3768 243051 3770
rect 150065 3712 150070 3768
rect 150126 3712 242990 3768
rect 243046 3712 243051 3768
rect 150065 3710 243051 3712
rect 150065 3707 150131 3710
rect 242985 3707 243051 3710
rect 140998 3572 141004 3636
rect 141068 3634 141074 3636
rect 148317 3634 148383 3637
rect 141068 3632 148383 3634
rect 141068 3576 148322 3632
rect 148378 3576 148383 3632
rect 141068 3574 148383 3576
rect 141068 3572 141074 3574
rect 148317 3571 148383 3574
rect 150525 3634 150591 3637
rect 264145 3634 264211 3637
rect 150525 3632 264211 3634
rect 150525 3576 150530 3632
rect 150586 3576 264150 3632
rect 264206 3576 264211 3632
rect 150525 3574 264211 3576
rect 150525 3571 150591 3574
rect 264145 3571 264211 3574
rect 143390 3436 143396 3500
rect 143460 3498 143466 3500
rect 164877 3498 164943 3501
rect 143460 3496 164943 3498
rect 143460 3440 164882 3496
rect 164938 3440 164943 3496
rect 143460 3438 164943 3440
rect 143460 3436 143466 3438
rect 164877 3435 164943 3438
rect 177062 3436 177068 3500
rect 177132 3498 177138 3500
rect 523033 3498 523099 3501
rect 177132 3496 523099 3498
rect 177132 3440 523038 3496
rect 523094 3440 523099 3496
rect 177132 3438 523099 3440
rect 177132 3436 177138 3438
rect 523033 3435 523099 3438
rect 101029 3362 101095 3365
rect 138054 3362 138060 3364
rect 101029 3360 138060 3362
rect 101029 3304 101034 3360
rect 101090 3304 138060 3360
rect 101029 3302 138060 3304
rect 101029 3299 101095 3302
rect 138054 3300 138060 3302
rect 138124 3300 138130 3364
rect 140814 3300 140820 3364
rect 140884 3362 140890 3364
rect 168373 3362 168439 3365
rect 140884 3360 168439 3362
rect 140884 3304 168378 3360
rect 168434 3304 168439 3360
rect 140884 3302 168439 3304
rect 140884 3300 140890 3302
rect 168373 3299 168439 3302
rect 176878 3300 176884 3364
rect 176948 3362 176954 3364
rect 562041 3362 562107 3365
rect 176948 3360 562107 3362
rect 176948 3304 562046 3360
rect 562102 3304 562107 3360
rect 176948 3302 562107 3304
rect 176948 3300 176954 3302
rect 562041 3299 562107 3302
<< via3 >>
rect 580212 697172 580276 697236
rect 580396 643996 580460 644060
rect 580396 82316 580460 82380
rect 164372 80412 164436 80476
rect 140820 80140 140884 80204
rect 134196 80004 134260 80068
rect 131252 79868 131316 79932
rect 131988 79868 132052 79932
rect 132356 79906 132360 79932
rect 132360 79906 132416 79932
rect 132416 79906 132420 79932
rect 132356 79868 132420 79906
rect 132908 79906 132912 79932
rect 132912 79906 132968 79932
rect 132968 79906 132972 79932
rect 132908 79868 132972 79906
rect 134380 79868 134444 79932
rect 133092 79732 133156 79796
rect 134196 79732 134260 79796
rect 143212 80004 143276 80068
rect 135300 79868 135364 79932
rect 136220 79868 136284 79932
rect 137692 79868 137756 79932
rect 137876 79868 137940 79932
rect 134932 79732 134996 79796
rect 135484 79732 135548 79796
rect 135852 79732 135916 79796
rect 138428 79732 138492 79796
rect 138980 79928 139044 79932
rect 138980 79872 138984 79928
rect 138984 79872 139040 79928
rect 139040 79872 139044 79928
rect 138980 79868 139044 79872
rect 139348 79868 139412 79932
rect 148364 80140 148428 80204
rect 139716 79732 139780 79796
rect 141372 79868 141436 79932
rect 142660 79928 142724 79932
rect 142660 79872 142664 79928
rect 142664 79872 142720 79928
rect 142720 79872 142724 79928
rect 142660 79868 142724 79872
rect 143948 79868 144012 79932
rect 144684 79928 144748 79932
rect 144684 79872 144688 79928
rect 144688 79872 144744 79928
rect 144744 79872 144748 79928
rect 144684 79868 144748 79872
rect 145236 79868 145300 79932
rect 146892 79868 146956 79932
rect 141004 79732 141068 79796
rect 143396 79792 143460 79796
rect 143396 79736 143446 79792
rect 143446 79736 143460 79792
rect 143396 79732 143460 79736
rect 144132 79732 144196 79796
rect 146524 79792 146588 79796
rect 146524 79736 146528 79792
rect 146528 79736 146584 79792
rect 146584 79736 146588 79792
rect 146524 79732 146588 79736
rect 147076 79732 147140 79796
rect 148180 79868 148244 79932
rect 151308 80140 151372 80204
rect 177988 80276 178052 80340
rect 149100 79906 149104 79932
rect 149104 79906 149160 79932
rect 149160 79906 149164 79932
rect 149100 79868 149164 79906
rect 149468 79868 149532 79932
rect 148732 79732 148796 79796
rect 149836 79732 149900 79796
rect 150756 79906 150760 79932
rect 150760 79906 150816 79932
rect 150816 79906 150820 79932
rect 150756 79868 150820 79906
rect 151124 79868 151188 79932
rect 151676 79906 151680 79932
rect 151680 79906 151736 79932
rect 151736 79906 151740 79932
rect 151676 79868 151740 79906
rect 152228 79868 152292 79932
rect 152964 79868 153028 79932
rect 153700 79928 153764 79932
rect 153700 79872 153704 79928
rect 153704 79872 153760 79928
rect 153760 79872 153764 79928
rect 153700 79868 153764 79872
rect 154068 79868 154132 79932
rect 154620 79868 154684 79932
rect 152412 79732 152476 79796
rect 155540 79906 155544 79932
rect 155544 79906 155600 79932
rect 155600 79906 155604 79932
rect 155540 79868 155604 79906
rect 155908 79868 155972 79932
rect 156460 79906 156464 79932
rect 156464 79906 156520 79932
rect 156520 79906 156524 79932
rect 156460 79868 156524 79906
rect 157012 79868 157076 79932
rect 156644 79792 156708 79796
rect 156644 79736 156648 79792
rect 156648 79736 156704 79792
rect 156704 79736 156708 79792
rect 156644 79732 156708 79736
rect 156828 79732 156892 79796
rect 168604 80140 168668 80204
rect 163820 80004 163884 80068
rect 171364 80004 171428 80068
rect 174308 80004 174372 80068
rect 157932 79906 157936 79932
rect 157936 79906 157992 79932
rect 157992 79906 157996 79932
rect 157932 79868 157996 79906
rect 158300 79868 158364 79932
rect 158116 79732 158180 79796
rect 158484 79596 158548 79660
rect 160508 79906 160512 79932
rect 160512 79906 160568 79932
rect 160568 79906 160572 79932
rect 160508 79868 160572 79906
rect 161244 79868 161308 79932
rect 161612 79928 161676 79932
rect 161612 79872 161616 79928
rect 161616 79872 161672 79928
rect 161672 79872 161676 79928
rect 161612 79868 161676 79872
rect 161980 79906 161984 79932
rect 161984 79906 162040 79932
rect 162040 79906 162044 79932
rect 161980 79868 162044 79906
rect 162348 79906 162352 79932
rect 162352 79906 162408 79932
rect 162408 79906 162412 79932
rect 162348 79868 162412 79906
rect 162716 79906 162720 79932
rect 162720 79906 162776 79932
rect 162776 79906 162780 79932
rect 162716 79868 162780 79906
rect 163636 79906 163640 79932
rect 163640 79906 163696 79932
rect 163696 79906 163700 79932
rect 163636 79868 163700 79906
rect 164372 79906 164376 79932
rect 164376 79906 164432 79932
rect 164432 79906 164436 79932
rect 164372 79868 164436 79906
rect 164004 79732 164068 79796
rect 164924 79868 164988 79932
rect 166580 79928 166644 79932
rect 166580 79872 166584 79928
rect 166584 79872 166640 79928
rect 166640 79872 166644 79928
rect 166580 79868 166644 79872
rect 166764 79868 166828 79932
rect 167316 79868 167380 79932
rect 162532 79596 162596 79660
rect 163084 79596 163148 79660
rect 164924 79596 164988 79660
rect 168052 79868 168116 79932
rect 169156 79928 169220 79932
rect 169156 79872 169160 79928
rect 169160 79872 169216 79928
rect 169216 79872 169220 79928
rect 169156 79868 169220 79872
rect 169524 79868 169588 79932
rect 170076 79906 170080 79932
rect 170080 79906 170136 79932
rect 170136 79906 170140 79932
rect 170076 79868 170140 79906
rect 172100 79868 172164 79932
rect 173388 79928 173452 79932
rect 173388 79872 173392 79928
rect 173392 79872 173448 79928
rect 173448 79872 173452 79928
rect 173388 79868 173452 79872
rect 173756 79906 173760 79932
rect 173760 79906 173816 79932
rect 173816 79906 173820 79932
rect 173756 79868 173820 79906
rect 174124 79906 174128 79932
rect 174128 79906 174184 79932
rect 174184 79906 174188 79932
rect 174124 79868 174188 79906
rect 174676 79928 174740 79932
rect 174676 79872 174680 79928
rect 174680 79872 174736 79928
rect 174736 79872 174740 79928
rect 174676 79868 174740 79872
rect 177068 80004 177132 80068
rect 175228 79906 175232 79932
rect 175232 79906 175288 79932
rect 175288 79906 175292 79932
rect 175228 79868 175292 79906
rect 170628 79732 170692 79796
rect 171548 79732 171612 79796
rect 174492 79732 174556 79796
rect 175780 79906 175784 79932
rect 175784 79906 175840 79932
rect 175840 79906 175844 79932
rect 175780 79868 175844 79906
rect 176332 79732 176396 79796
rect 178540 79928 178604 79932
rect 178540 79872 178544 79928
rect 178544 79872 178600 79928
rect 178600 79872 178604 79928
rect 166396 79596 166460 79660
rect 166764 79596 166828 79660
rect 167868 79596 167932 79660
rect 178540 79868 178604 79872
rect 177988 79656 178052 79660
rect 177988 79600 178038 79656
rect 178038 79600 178052 79656
rect 177988 79596 178052 79600
rect 168604 79520 168668 79524
rect 168604 79464 168618 79520
rect 168618 79464 168668 79520
rect 168604 79460 168668 79464
rect 170444 79520 170508 79524
rect 170444 79464 170494 79520
rect 170494 79464 170508 79520
rect 170444 79460 170508 79464
rect 171916 79460 171980 79524
rect 173388 79520 173452 79524
rect 173388 79464 173402 79520
rect 173402 79464 173452 79520
rect 173388 79460 173452 79464
rect 580212 79324 580276 79388
rect 155540 79052 155604 79116
rect 162164 79052 162228 79116
rect 163636 79052 163700 79116
rect 138980 78916 139044 78980
rect 156644 78976 156708 78980
rect 156644 78920 156694 78976
rect 156694 78920 156708 78976
rect 156644 78916 156708 78920
rect 158852 78916 158916 78980
rect 162348 78976 162412 78980
rect 162348 78920 162362 78976
rect 162362 78920 162412 78976
rect 162348 78916 162412 78920
rect 164004 78976 164068 78980
rect 164004 78920 164054 78976
rect 164054 78920 164068 78976
rect 164004 78916 164068 78920
rect 136588 78780 136652 78844
rect 138060 78780 138124 78844
rect 160692 78780 160756 78844
rect 161980 78840 162044 78844
rect 161980 78784 161994 78840
rect 161994 78784 162044 78840
rect 134932 78644 134996 78708
rect 136220 78704 136284 78708
rect 136220 78648 136234 78704
rect 136234 78648 136284 78704
rect 136220 78644 136284 78648
rect 137508 78644 137572 78708
rect 137692 78704 137756 78708
rect 137692 78648 137742 78704
rect 137742 78648 137756 78704
rect 137692 78644 137756 78648
rect 138244 78644 138308 78708
rect 139532 78704 139596 78708
rect 139532 78648 139546 78704
rect 139546 78648 139596 78704
rect 139532 78644 139596 78648
rect 141372 78644 141436 78708
rect 160876 78644 160940 78708
rect 161980 78780 162044 78784
rect 163268 78780 163332 78844
rect 166580 78780 166644 78844
rect 166764 78840 166828 78844
rect 167684 78916 167748 78980
rect 174860 79052 174924 79116
rect 178540 79188 178604 79252
rect 166764 78784 166778 78840
rect 166778 78784 166828 78840
rect 166764 78780 166828 78784
rect 161612 78644 161676 78708
rect 162348 78644 162412 78708
rect 163084 78644 163148 78708
rect 163452 78644 163516 78708
rect 165108 78644 165172 78708
rect 165476 78704 165540 78708
rect 165476 78648 165526 78704
rect 165526 78648 165540 78704
rect 165476 78644 165540 78648
rect 166580 78644 166644 78708
rect 167500 78644 167564 78708
rect 169708 78704 169772 78708
rect 169708 78648 169722 78704
rect 169722 78648 169772 78704
rect 169708 78644 169772 78648
rect 170996 78704 171060 78708
rect 170996 78648 171046 78704
rect 171046 78648 171060 78704
rect 170996 78644 171060 78648
rect 171732 78644 171796 78708
rect 175228 78704 175292 78708
rect 175228 78648 175242 78704
rect 175242 78648 175292 78704
rect 175228 78644 175292 78648
rect 175964 78704 176028 78708
rect 175964 78648 176014 78704
rect 176014 78648 176028 78704
rect 175964 78644 176028 78648
rect 150756 78236 150820 78300
rect 166212 78236 166276 78300
rect 172100 78568 172164 78572
rect 172100 78512 172150 78568
rect 172150 78512 172164 78568
rect 172100 78508 172164 78512
rect 172100 78372 172164 78436
rect 174676 78372 174740 78436
rect 176516 78372 176580 78436
rect 132356 78100 132420 78164
rect 132908 78160 132972 78164
rect 132908 78104 132922 78160
rect 132922 78104 132972 78160
rect 132908 78100 132972 78104
rect 139164 78100 139228 78164
rect 167316 78100 167380 78164
rect 174308 78100 174372 78164
rect 174676 78100 174740 78164
rect 131988 77828 132052 77892
rect 137876 77828 137940 77892
rect 170260 77828 170324 77892
rect 174124 77888 174188 77892
rect 174124 77832 174174 77888
rect 174174 77832 174188 77888
rect 174124 77828 174188 77832
rect 176884 77828 176948 77892
rect 141004 77556 141068 77620
rect 144500 77556 144564 77620
rect 142844 77420 142908 77484
rect 144316 77420 144380 77484
rect 145236 77420 145300 77484
rect 145420 77420 145484 77484
rect 147444 77480 147508 77484
rect 147444 77424 147494 77480
rect 147494 77424 147508 77480
rect 135484 77344 135548 77348
rect 135484 77288 135534 77344
rect 135534 77288 135548 77344
rect 135484 77284 135548 77288
rect 140636 77284 140700 77348
rect 131620 77148 131684 77212
rect 143028 77284 143092 77348
rect 145236 77284 145300 77348
rect 147444 77420 147508 77424
rect 146892 77284 146956 77348
rect 147260 77284 147324 77348
rect 161244 77344 161308 77348
rect 161244 77288 161294 77344
rect 161294 77288 161308 77344
rect 161244 77284 161308 77288
rect 173572 77284 173636 77348
rect 177068 77556 177132 77620
rect 170444 77208 170508 77212
rect 170444 77152 170458 77208
rect 170458 77152 170508 77208
rect 170444 77148 170508 77152
rect 153884 77012 153948 77076
rect 157932 76876 157996 76940
rect 160508 76876 160572 76940
rect 145604 76740 145668 76804
rect 141004 76604 141068 76668
rect 142660 76604 142724 76668
rect 143948 76604 144012 76668
rect 146524 76604 146588 76668
rect 148180 76604 148244 76668
rect 149652 76604 149716 76668
rect 139348 76468 139412 76532
rect 156828 76196 156892 76260
rect 148916 76060 148980 76124
rect 149468 76120 149532 76124
rect 149468 76064 149482 76120
rect 149482 76064 149532 76120
rect 149468 76060 149532 76064
rect 152780 76060 152844 76124
rect 156644 76060 156708 76124
rect 171364 76060 171428 76124
rect 177068 76060 177132 76124
rect 148548 75924 148612 75988
rect 149100 75924 149164 75988
rect 150020 75984 150084 75988
rect 150020 75928 150034 75984
rect 150034 75928 150084 75984
rect 150020 75924 150084 75928
rect 151124 75924 151188 75988
rect 151492 75924 151556 75988
rect 152228 75984 152292 75988
rect 152228 75928 152242 75984
rect 152242 75928 152292 75984
rect 152228 75924 152292 75928
rect 152964 75924 153028 75988
rect 153700 75924 153764 75988
rect 154252 75924 154316 75988
rect 154620 75924 154684 75988
rect 169156 75924 169220 75988
rect 170076 75924 170140 75988
rect 170812 75984 170876 75988
rect 170812 75928 170862 75984
rect 170862 75928 170876 75984
rect 170812 75924 170876 75928
rect 171548 75924 171612 75988
rect 175964 75924 176028 75988
rect 133276 75788 133340 75852
rect 144684 75788 144748 75852
rect 136588 75380 136652 75444
rect 155908 74972 155972 75036
rect 160876 74564 160940 74628
rect 161428 74564 161492 74628
rect 157012 74292 157076 74356
rect 161244 74156 161308 74220
rect 135852 73748 135916 73812
rect 156460 73748 156524 73812
rect 174492 73476 174556 73540
rect 131068 73264 131132 73268
rect 131068 73208 131118 73264
rect 131118 73208 131132 73264
rect 131068 73204 131132 73208
rect 138428 72660 138492 72724
rect 158300 72524 158364 72588
rect 131620 72388 131684 72452
rect 168052 72388 168116 72452
rect 158116 71708 158180 71772
rect 156644 71572 156708 71636
rect 158852 71436 158916 71500
rect 161428 71300 161492 71364
rect 169708 71164 169772 71228
rect 170628 71028 170692 71092
rect 167684 69532 167748 69596
rect 144316 68444 144380 68508
rect 158484 68308 158548 68372
rect 167868 68172 167932 68236
rect 144500 66812 144564 66876
rect 145236 63004 145300 63068
rect 174860 62868 174924 62932
rect 176148 62732 176212 62796
rect 171916 61508 171980 61572
rect 176332 61372 176396 61436
rect 144132 57156 144196 57220
rect 161060 48860 161124 48924
rect 176516 46140 176580 46204
rect 131252 35124 131316 35188
rect 147076 34172 147140 34236
rect 163452 34036 163516 34100
rect 163268 33900 163332 33964
rect 173572 33764 173636 33828
rect 163636 31316 163700 31380
rect 166212 31180 166276 31244
rect 167500 31044 167564 31108
rect 173756 30908 173820 30972
rect 151308 28460 151372 28524
rect 166396 28324 166460 28388
rect 145420 25468 145484 25532
rect 170812 24244 170876 24308
rect 174676 24108 174740 24172
rect 147260 23292 147324 23356
rect 152412 23156 152476 23220
rect 140636 23020 140700 23084
rect 170260 22884 170324 22948
rect 170996 22748 171060 22812
rect 135668 22612 135732 22676
rect 172100 22612 172164 22676
rect 169524 21252 169588 21316
rect 145604 20436 145668 20500
rect 139164 20300 139228 20364
rect 162348 20164 162412 20228
rect 162164 20028 162228 20092
rect 171732 19892 171796 19956
rect 142844 18668 142908 18732
rect 148364 18532 148428 18596
rect 165292 17716 165356 17780
rect 165108 17580 165172 17644
rect 164924 17444 164988 17508
rect 166764 17308 166828 17372
rect 166580 17172 166644 17236
rect 152596 14452 152660 14516
rect 149652 12004 149716 12068
rect 151492 11868 151556 11932
rect 162532 11732 162596 11796
rect 139532 11596 139596 11660
rect 162716 11596 162780 11660
rect 138244 10372 138308 10436
rect 148548 10372 148612 10436
rect 137508 10236 137572 10300
rect 160692 10236 160756 10300
rect 153884 9148 153948 9212
rect 139716 9012 139780 9076
rect 154068 9012 154132 9076
rect 134196 8876 134260 8940
rect 154252 8876 154316 8940
rect 135484 7924 135548 7988
rect 135300 7788 135364 7852
rect 134012 7652 134076 7716
rect 134380 7516 134444 7580
rect 150020 6836 150084 6900
rect 149836 6700 149900 6764
rect 151676 6564 151740 6628
rect 131068 6428 131132 6492
rect 152964 6428 153028 6492
rect 133092 6292 133156 6356
rect 152780 6292 152844 6356
rect 133276 6156 133340 6220
rect 165476 6156 165540 6220
rect 147444 6020 147508 6084
rect 143028 4932 143092 4996
rect 143212 4796 143276 4860
rect 148732 3980 148796 4044
rect 148916 3844 148980 3908
rect 141004 3572 141068 3636
rect 143396 3436 143460 3500
rect 177068 3436 177132 3500
rect 138060 3300 138124 3364
rect 140820 3300 140884 3364
rect 176884 3300 176948 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 628954 51914 664398
rect 51294 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 51914 628954
rect 51294 628634 51914 628718
rect 51294 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 51914 628634
rect 51294 592954 51914 628398
rect 51294 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 51914 592954
rect 51294 592634 51914 592718
rect 51294 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 51914 592634
rect 51294 556954 51914 592398
rect 51294 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 51914 556954
rect 51294 556634 51914 556718
rect 51294 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 51914 556634
rect 51294 520954 51914 556398
rect 51294 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 51914 520954
rect 51294 520634 51914 520718
rect 51294 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 51914 520634
rect 51294 484954 51914 520398
rect 51294 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 51914 484954
rect 51294 484634 51914 484718
rect 51294 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 51914 484634
rect 51294 448954 51914 484398
rect 51294 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 51914 448954
rect 51294 448634 51914 448718
rect 51294 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 51914 448634
rect 51294 412954 51914 448398
rect 51294 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 51914 412954
rect 51294 412634 51914 412718
rect 51294 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 51914 412634
rect 51294 376954 51914 412398
rect 51294 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 51914 376954
rect 51294 376634 51914 376718
rect 51294 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 51914 376634
rect 51294 340954 51914 376398
rect 51294 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 51914 340954
rect 51294 340634 51914 340718
rect 51294 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 51914 340634
rect 51294 304954 51914 340398
rect 51294 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 51914 304954
rect 51294 304634 51914 304718
rect 51294 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 51914 304634
rect 51294 268954 51914 304398
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 51294 196954 51914 232398
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 637954 60914 673398
rect 60294 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 60914 637954
rect 60294 637634 60914 637718
rect 60294 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 60914 637634
rect 60294 601954 60914 637398
rect 60294 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 60914 601954
rect 60294 601634 60914 601718
rect 60294 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 60914 601634
rect 60294 565954 60914 601398
rect 60294 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 60914 565954
rect 60294 565634 60914 565718
rect 60294 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 60914 565634
rect 60294 529954 60914 565398
rect 60294 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 60914 529954
rect 60294 529634 60914 529718
rect 60294 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 60914 529634
rect 60294 493954 60914 529398
rect 60294 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 60914 493954
rect 60294 493634 60914 493718
rect 60294 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 60914 493634
rect 60294 457954 60914 493398
rect 60294 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 60914 457954
rect 60294 457634 60914 457718
rect 60294 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 60914 457634
rect 60294 421954 60914 457398
rect 60294 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 60914 421954
rect 60294 421634 60914 421718
rect 60294 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 60914 421634
rect 60294 385954 60914 421398
rect 60294 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 60914 385954
rect 60294 385634 60914 385718
rect 60294 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 60914 385634
rect 60294 349954 60914 385398
rect 60294 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 60914 349954
rect 60294 349634 60914 349718
rect 60294 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 60914 349634
rect 60294 313954 60914 349398
rect 60294 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 60914 313954
rect 60294 313634 60914 313718
rect 60294 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 60914 313634
rect 60294 277954 60914 313398
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 60294 205954 60914 241398
rect 60294 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 60914 205954
rect 60294 205634 60914 205718
rect 60294 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 60914 205634
rect 60294 169954 60914 205398
rect 60294 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 60914 169954
rect 60294 169634 60914 169718
rect 60294 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 60914 169634
rect 60294 133954 60914 169398
rect 60294 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 60914 133954
rect 60294 133634 60914 133718
rect 60294 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 60914 133634
rect 60294 97954 60914 133398
rect 60294 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 60914 97954
rect 60294 97634 60914 97718
rect 60294 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 60914 97634
rect 60294 61954 60914 97398
rect 60294 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 60914 61954
rect 60294 61634 60914 61718
rect 60294 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 60914 61634
rect 60294 25954 60914 61398
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 642454 65414 677898
rect 64794 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 65414 642454
rect 64794 642134 65414 642218
rect 64794 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 65414 642134
rect 64794 606454 65414 641898
rect 64794 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 65414 606454
rect 64794 606134 65414 606218
rect 64794 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 65414 606134
rect 64794 570454 65414 605898
rect 64794 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 65414 570454
rect 64794 570134 65414 570218
rect 64794 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 65414 570134
rect 64794 534454 65414 569898
rect 64794 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 65414 534454
rect 64794 534134 65414 534218
rect 64794 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 65414 534134
rect 64794 498454 65414 533898
rect 64794 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 65414 498454
rect 64794 498134 65414 498218
rect 64794 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 65414 498134
rect 64794 462454 65414 497898
rect 64794 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 65414 462454
rect 64794 462134 65414 462218
rect 64794 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 65414 462134
rect 64794 426454 65414 461898
rect 64794 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 65414 426454
rect 64794 426134 65414 426218
rect 64794 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 65414 426134
rect 64794 390454 65414 425898
rect 64794 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 65414 390454
rect 64794 390134 65414 390218
rect 64794 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 65414 390134
rect 64794 354454 65414 389898
rect 64794 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 65414 354454
rect 64794 354134 65414 354218
rect 64794 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 65414 354134
rect 64794 318454 65414 353898
rect 64794 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 65414 318454
rect 64794 318134 65414 318218
rect 64794 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 65414 318134
rect 64794 282454 65414 317898
rect 64794 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 65414 282454
rect 64794 282134 65414 282218
rect 64794 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 65414 282134
rect 64794 246454 65414 281898
rect 64794 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 65414 246454
rect 64794 246134 65414 246218
rect 64794 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 65414 246134
rect 64794 210454 65414 245898
rect 64794 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 65414 210454
rect 64794 210134 65414 210218
rect 64794 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 65414 210134
rect 64794 174454 65414 209898
rect 64794 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 65414 174454
rect 64794 174134 65414 174218
rect 64794 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 65414 174134
rect 64794 138454 65414 173898
rect 64794 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 65414 138454
rect 64794 138134 65414 138218
rect 64794 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 65414 138134
rect 64794 102454 65414 137898
rect 64794 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 65414 102454
rect 64794 102134 65414 102218
rect 64794 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 65414 102134
rect 64794 66454 65414 101898
rect 64794 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 65414 66454
rect 64794 66134 65414 66218
rect 64794 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 65414 66134
rect 64794 30454 65414 65898
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 646954 69914 682398
rect 69294 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 69914 646954
rect 69294 646634 69914 646718
rect 69294 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 69914 646634
rect 69294 610954 69914 646398
rect 69294 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 69914 610954
rect 69294 610634 69914 610718
rect 69294 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 69914 610634
rect 69294 574954 69914 610398
rect 69294 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 69914 574954
rect 69294 574634 69914 574718
rect 69294 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 69914 574634
rect 69294 538954 69914 574398
rect 69294 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 69914 538954
rect 69294 538634 69914 538718
rect 69294 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 69914 538634
rect 69294 502954 69914 538398
rect 69294 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 69914 502954
rect 69294 502634 69914 502718
rect 69294 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 69914 502634
rect 69294 466954 69914 502398
rect 69294 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 69914 466954
rect 69294 466634 69914 466718
rect 69294 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 69914 466634
rect 69294 430954 69914 466398
rect 69294 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 69914 430954
rect 69294 430634 69914 430718
rect 69294 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 69914 430634
rect 69294 394954 69914 430398
rect 69294 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 69914 394954
rect 69294 394634 69914 394718
rect 69294 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 69914 394634
rect 69294 358954 69914 394398
rect 69294 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 69914 358954
rect 69294 358634 69914 358718
rect 69294 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 69914 358634
rect 69294 322954 69914 358398
rect 69294 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 69914 322954
rect 69294 322634 69914 322718
rect 69294 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 69914 322634
rect 69294 286954 69914 322398
rect 69294 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 69914 286954
rect 69294 286634 69914 286718
rect 69294 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 69914 286634
rect 69294 250954 69914 286398
rect 69294 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 69914 250954
rect 69294 250634 69914 250718
rect 69294 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 69914 250634
rect 69294 214954 69914 250398
rect 69294 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 69914 214954
rect 69294 214634 69914 214718
rect 69294 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 69914 214634
rect 69294 178954 69914 214398
rect 69294 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 69914 178954
rect 69294 178634 69914 178718
rect 69294 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 69914 178634
rect 69294 142954 69914 178398
rect 69294 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 69914 142954
rect 69294 142634 69914 142718
rect 69294 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 69914 142634
rect 69294 106954 69914 142398
rect 69294 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 69914 106954
rect 69294 106634 69914 106718
rect 69294 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 69914 106634
rect 69294 70954 69914 106398
rect 69294 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 69914 70954
rect 69294 70634 69914 70718
rect 69294 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 69914 70634
rect 69294 34954 69914 70398
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 655954 78914 691398
rect 78294 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 78914 655954
rect 78294 655634 78914 655718
rect 78294 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 78914 655634
rect 78294 619954 78914 655398
rect 78294 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 78914 619954
rect 78294 619634 78914 619718
rect 78294 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 78914 619634
rect 78294 583954 78914 619398
rect 78294 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 78914 583954
rect 78294 583634 78914 583718
rect 78294 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 78914 583634
rect 78294 547954 78914 583398
rect 78294 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 78914 547954
rect 78294 547634 78914 547718
rect 78294 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 78914 547634
rect 78294 511954 78914 547398
rect 78294 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 78914 511954
rect 78294 511634 78914 511718
rect 78294 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 78914 511634
rect 78294 475954 78914 511398
rect 78294 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 78914 475954
rect 78294 475634 78914 475718
rect 78294 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 78914 475634
rect 78294 439954 78914 475398
rect 78294 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 78914 439954
rect 78294 439634 78914 439718
rect 78294 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 78914 439634
rect 78294 403954 78914 439398
rect 78294 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 78914 403954
rect 78294 403634 78914 403718
rect 78294 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 78914 403634
rect 78294 367954 78914 403398
rect 78294 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 78914 367954
rect 78294 367634 78914 367718
rect 78294 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 78914 367634
rect 78294 331954 78914 367398
rect 78294 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 78914 331954
rect 78294 331634 78914 331718
rect 78294 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 78914 331634
rect 78294 295954 78914 331398
rect 78294 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 78914 295954
rect 78294 295634 78914 295718
rect 78294 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 78914 295634
rect 78294 259954 78914 295398
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 187954 78914 223398
rect 78294 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 78914 187954
rect 78294 187634 78914 187718
rect 78294 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 78914 187634
rect 78294 151954 78914 187398
rect 78294 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 78914 151954
rect 78294 151634 78914 151718
rect 78294 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 78914 151634
rect 78294 115954 78914 151398
rect 78294 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 78914 115954
rect 78294 115634 78914 115718
rect 78294 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 78914 115634
rect 78294 79954 78914 115398
rect 78294 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 78914 79954
rect 78294 79634 78914 79718
rect 78294 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 78914 79634
rect 78294 43954 78914 79398
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 660454 83414 695898
rect 82794 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 83414 660454
rect 82794 660134 83414 660218
rect 82794 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 83414 660134
rect 82794 624454 83414 659898
rect 82794 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 83414 624454
rect 82794 624134 83414 624218
rect 82794 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 83414 624134
rect 82794 588454 83414 623898
rect 82794 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 83414 588454
rect 82794 588134 83414 588218
rect 82794 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 83414 588134
rect 82794 552454 83414 587898
rect 82794 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 83414 552454
rect 82794 552134 83414 552218
rect 82794 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 83414 552134
rect 82794 516454 83414 551898
rect 82794 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 83414 516454
rect 82794 516134 83414 516218
rect 82794 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 83414 516134
rect 82794 480454 83414 515898
rect 82794 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 83414 480454
rect 82794 480134 83414 480218
rect 82794 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 83414 480134
rect 82794 444454 83414 479898
rect 82794 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 83414 444454
rect 82794 444134 83414 444218
rect 82794 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 83414 444134
rect 82794 408454 83414 443898
rect 82794 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 83414 408454
rect 82794 408134 83414 408218
rect 82794 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 83414 408134
rect 82794 372454 83414 407898
rect 82794 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 83414 372454
rect 82794 372134 83414 372218
rect 82794 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 83414 372134
rect 82794 336454 83414 371898
rect 82794 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 83414 336454
rect 82794 336134 83414 336218
rect 82794 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 83414 336134
rect 82794 300454 83414 335898
rect 82794 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 83414 300454
rect 82794 300134 83414 300218
rect 82794 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 83414 300134
rect 82794 264454 83414 299898
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 192454 83414 227898
rect 82794 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 83414 192454
rect 82794 192134 83414 192218
rect 82794 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 83414 192134
rect 82794 156454 83414 191898
rect 82794 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 83414 156454
rect 82794 156134 83414 156218
rect 82794 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 83414 156134
rect 82794 120454 83414 155898
rect 82794 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 83414 120454
rect 82794 120134 83414 120218
rect 82794 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 83414 120134
rect 82794 84454 83414 119898
rect 82794 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 83414 84454
rect 82794 84134 83414 84218
rect 82794 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 83414 84134
rect 82794 48454 83414 83898
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 628954 87914 664398
rect 87294 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 87914 628954
rect 87294 628634 87914 628718
rect 87294 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 87914 628634
rect 87294 592954 87914 628398
rect 87294 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 87914 592954
rect 87294 592634 87914 592718
rect 87294 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 87914 592634
rect 87294 556954 87914 592398
rect 87294 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 87914 556954
rect 87294 556634 87914 556718
rect 87294 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 87914 556634
rect 87294 520954 87914 556398
rect 87294 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 87914 520954
rect 87294 520634 87914 520718
rect 87294 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 87914 520634
rect 87294 484954 87914 520398
rect 87294 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 87914 484954
rect 87294 484634 87914 484718
rect 87294 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 87914 484634
rect 87294 448954 87914 484398
rect 87294 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 87914 448954
rect 87294 448634 87914 448718
rect 87294 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 87914 448634
rect 87294 412954 87914 448398
rect 87294 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 87914 412954
rect 87294 412634 87914 412718
rect 87294 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 87914 412634
rect 87294 376954 87914 412398
rect 87294 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 87914 376954
rect 87294 376634 87914 376718
rect 87294 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 87914 376634
rect 87294 340954 87914 376398
rect 87294 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 87914 340954
rect 87294 340634 87914 340718
rect 87294 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 87914 340634
rect 87294 304954 87914 340398
rect 87294 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 87914 304954
rect 87294 304634 87914 304718
rect 87294 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 87914 304634
rect 87294 268954 87914 304398
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 196954 87914 232398
rect 87294 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 87914 196954
rect 87294 196634 87914 196718
rect 87294 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 87914 196634
rect 87294 160954 87914 196398
rect 87294 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 87914 160954
rect 87294 160634 87914 160718
rect 87294 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 87914 160634
rect 87294 124954 87914 160398
rect 87294 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 87914 124954
rect 87294 124634 87914 124718
rect 87294 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 87914 124634
rect 87294 88954 87914 124398
rect 87294 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 87914 88954
rect 87294 88634 87914 88718
rect 87294 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 87914 88634
rect 87294 52954 87914 88398
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 637954 96914 673398
rect 96294 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 96914 637954
rect 96294 637634 96914 637718
rect 96294 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 96914 637634
rect 96294 601954 96914 637398
rect 96294 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 96914 601954
rect 96294 601634 96914 601718
rect 96294 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 96914 601634
rect 96294 565954 96914 601398
rect 96294 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 96914 565954
rect 96294 565634 96914 565718
rect 96294 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 96914 565634
rect 96294 529954 96914 565398
rect 96294 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 96914 529954
rect 96294 529634 96914 529718
rect 96294 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 96914 529634
rect 96294 493954 96914 529398
rect 96294 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 96914 493954
rect 96294 493634 96914 493718
rect 96294 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 96914 493634
rect 96294 457954 96914 493398
rect 96294 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 96914 457954
rect 96294 457634 96914 457718
rect 96294 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 96914 457634
rect 96294 421954 96914 457398
rect 96294 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 96914 421954
rect 96294 421634 96914 421718
rect 96294 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 96914 421634
rect 96294 385954 96914 421398
rect 96294 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 96914 385954
rect 96294 385634 96914 385718
rect 96294 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 96914 385634
rect 96294 349954 96914 385398
rect 96294 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 96914 349954
rect 96294 349634 96914 349718
rect 96294 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 96914 349634
rect 96294 313954 96914 349398
rect 96294 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 96914 313954
rect 96294 313634 96914 313718
rect 96294 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 96914 313634
rect 96294 277954 96914 313398
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 205954 96914 241398
rect 96294 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 96914 205954
rect 96294 205634 96914 205718
rect 96294 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 96914 205634
rect 96294 169954 96914 205398
rect 96294 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 96914 169954
rect 96294 169634 96914 169718
rect 96294 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 96914 169634
rect 96294 133954 96914 169398
rect 96294 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 96914 133954
rect 96294 133634 96914 133718
rect 96294 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 96914 133634
rect 96294 97954 96914 133398
rect 96294 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 96914 97954
rect 96294 97634 96914 97718
rect 96294 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 96914 97634
rect 96294 61954 96914 97398
rect 96294 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 96914 61954
rect 96294 61634 96914 61718
rect 96294 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 96914 61634
rect 96294 25954 96914 61398
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 642454 101414 677898
rect 100794 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 101414 642454
rect 100794 642134 101414 642218
rect 100794 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 101414 642134
rect 100794 606454 101414 641898
rect 100794 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 101414 606454
rect 100794 606134 101414 606218
rect 100794 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 101414 606134
rect 100794 570454 101414 605898
rect 100794 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 101414 570454
rect 100794 570134 101414 570218
rect 100794 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 101414 570134
rect 100794 534454 101414 569898
rect 100794 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 101414 534454
rect 100794 534134 101414 534218
rect 100794 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 101414 534134
rect 100794 498454 101414 533898
rect 100794 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 101414 498454
rect 100794 498134 101414 498218
rect 100794 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 101414 498134
rect 100794 462454 101414 497898
rect 100794 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 101414 462454
rect 100794 462134 101414 462218
rect 100794 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 101414 462134
rect 100794 426454 101414 461898
rect 100794 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 101414 426454
rect 100794 426134 101414 426218
rect 100794 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 101414 426134
rect 100794 390454 101414 425898
rect 100794 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 101414 390454
rect 100794 390134 101414 390218
rect 100794 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 101414 390134
rect 100794 354454 101414 389898
rect 100794 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 101414 354454
rect 100794 354134 101414 354218
rect 100794 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 101414 354134
rect 100794 318454 101414 353898
rect 100794 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 101414 318454
rect 100794 318134 101414 318218
rect 100794 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 101414 318134
rect 100794 282454 101414 317898
rect 100794 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 101414 282454
rect 100794 282134 101414 282218
rect 100794 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 101414 282134
rect 100794 246454 101414 281898
rect 100794 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 101414 246454
rect 100794 246134 101414 246218
rect 100794 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 101414 246134
rect 100794 210454 101414 245898
rect 100794 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 101414 210454
rect 100794 210134 101414 210218
rect 100794 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 101414 210134
rect 100794 174454 101414 209898
rect 100794 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 101414 174454
rect 100794 174134 101414 174218
rect 100794 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 101414 174134
rect 100794 138454 101414 173898
rect 100794 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 101414 138454
rect 100794 138134 101414 138218
rect 100794 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 101414 138134
rect 100794 102454 101414 137898
rect 100794 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 101414 102454
rect 100794 102134 101414 102218
rect 100794 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 101414 102134
rect 100794 66454 101414 101898
rect 100794 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 101414 66454
rect 100794 66134 101414 66218
rect 100794 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 101414 66134
rect 100794 30454 101414 65898
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 646954 105914 682398
rect 105294 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 105914 646954
rect 105294 646634 105914 646718
rect 105294 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 105914 646634
rect 105294 610954 105914 646398
rect 105294 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 105914 610954
rect 105294 610634 105914 610718
rect 105294 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 105914 610634
rect 105294 574954 105914 610398
rect 105294 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 105914 574954
rect 105294 574634 105914 574718
rect 105294 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 105914 574634
rect 105294 538954 105914 574398
rect 105294 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 105914 538954
rect 105294 538634 105914 538718
rect 105294 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 105914 538634
rect 105294 502954 105914 538398
rect 105294 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 105914 502954
rect 105294 502634 105914 502718
rect 105294 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 105914 502634
rect 105294 466954 105914 502398
rect 105294 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 105914 466954
rect 105294 466634 105914 466718
rect 105294 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 105914 466634
rect 105294 430954 105914 466398
rect 105294 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 105914 430954
rect 105294 430634 105914 430718
rect 105294 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 105914 430634
rect 105294 394954 105914 430398
rect 105294 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 105914 394954
rect 105294 394634 105914 394718
rect 105294 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 105914 394634
rect 105294 358954 105914 394398
rect 105294 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 105914 358954
rect 105294 358634 105914 358718
rect 105294 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 105914 358634
rect 105294 322954 105914 358398
rect 105294 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 105914 322954
rect 105294 322634 105914 322718
rect 105294 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 105914 322634
rect 105294 286954 105914 322398
rect 105294 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 105914 286954
rect 105294 286634 105914 286718
rect 105294 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 105914 286634
rect 105294 250954 105914 286398
rect 105294 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 105914 250954
rect 105294 250634 105914 250718
rect 105294 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 105914 250634
rect 105294 214954 105914 250398
rect 105294 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 105914 214954
rect 105294 214634 105914 214718
rect 105294 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 105914 214634
rect 105294 178954 105914 214398
rect 105294 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 105914 178954
rect 105294 178634 105914 178718
rect 105294 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 105914 178634
rect 105294 142954 105914 178398
rect 105294 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 105914 142954
rect 105294 142634 105914 142718
rect 105294 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 105914 142634
rect 105294 106954 105914 142398
rect 105294 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 105914 106954
rect 105294 106634 105914 106718
rect 105294 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 105914 106634
rect 105294 70954 105914 106398
rect 105294 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 105914 70954
rect 105294 70634 105914 70718
rect 105294 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 105914 70634
rect 105294 34954 105914 70398
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 655954 114914 691398
rect 114294 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 114914 655954
rect 114294 655634 114914 655718
rect 114294 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 114914 655634
rect 114294 619954 114914 655398
rect 114294 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 114914 619954
rect 114294 619634 114914 619718
rect 114294 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 114914 619634
rect 114294 583954 114914 619398
rect 114294 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 114914 583954
rect 114294 583634 114914 583718
rect 114294 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 114914 583634
rect 114294 547954 114914 583398
rect 114294 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 114914 547954
rect 114294 547634 114914 547718
rect 114294 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 114914 547634
rect 114294 511954 114914 547398
rect 114294 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 114914 511954
rect 114294 511634 114914 511718
rect 114294 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 114914 511634
rect 114294 475954 114914 511398
rect 114294 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 114914 475954
rect 114294 475634 114914 475718
rect 114294 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 114914 475634
rect 114294 439954 114914 475398
rect 114294 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 114914 439954
rect 114294 439634 114914 439718
rect 114294 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 114914 439634
rect 114294 403954 114914 439398
rect 114294 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 114914 403954
rect 114294 403634 114914 403718
rect 114294 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 114914 403634
rect 114294 367954 114914 403398
rect 114294 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 114914 367954
rect 114294 367634 114914 367718
rect 114294 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 114914 367634
rect 114294 331954 114914 367398
rect 114294 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 114914 331954
rect 114294 331634 114914 331718
rect 114294 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 114914 331634
rect 114294 295954 114914 331398
rect 114294 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 114914 295954
rect 114294 295634 114914 295718
rect 114294 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 114914 295634
rect 114294 259954 114914 295398
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 187954 114914 223398
rect 114294 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 114914 187954
rect 114294 187634 114914 187718
rect 114294 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 114914 187634
rect 114294 151954 114914 187398
rect 114294 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 114914 151954
rect 114294 151634 114914 151718
rect 114294 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 114914 151634
rect 114294 115954 114914 151398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 660454 119414 695898
rect 118794 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 119414 660454
rect 118794 660134 119414 660218
rect 118794 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 119414 660134
rect 118794 624454 119414 659898
rect 118794 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 119414 624454
rect 118794 624134 119414 624218
rect 118794 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 119414 624134
rect 118794 588454 119414 623898
rect 118794 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 119414 588454
rect 118794 588134 119414 588218
rect 118794 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 119414 588134
rect 118794 552454 119414 587898
rect 118794 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 119414 552454
rect 118794 552134 119414 552218
rect 118794 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 119414 552134
rect 118794 516454 119414 551898
rect 118794 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 119414 516454
rect 118794 516134 119414 516218
rect 118794 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 119414 516134
rect 118794 480454 119414 515898
rect 118794 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 119414 480454
rect 118794 480134 119414 480218
rect 118794 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 119414 480134
rect 118794 444454 119414 479898
rect 118794 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 119414 444454
rect 118794 444134 119414 444218
rect 118794 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 119414 444134
rect 118794 408454 119414 443898
rect 118794 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 119414 408454
rect 118794 408134 119414 408218
rect 118794 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 119414 408134
rect 118794 372454 119414 407898
rect 118794 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 119414 372454
rect 118794 372134 119414 372218
rect 118794 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 119414 372134
rect 118794 336454 119414 371898
rect 118794 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 119414 336454
rect 118794 336134 119414 336218
rect 118794 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 119414 336134
rect 118794 300454 119414 335898
rect 118794 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 119414 300454
rect 118794 300134 119414 300218
rect 118794 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 119414 300134
rect 118794 264454 119414 299898
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 192454 119414 227898
rect 118794 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 119414 192454
rect 118794 192134 119414 192218
rect 118794 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 119414 192134
rect 118794 156454 119414 191898
rect 118794 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 119414 156454
rect 118794 156134 119414 156218
rect 118794 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 119414 156134
rect 118794 142000 119414 155898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 628954 123914 664398
rect 123294 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 123914 628954
rect 123294 628634 123914 628718
rect 123294 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 123914 628634
rect 123294 592954 123914 628398
rect 123294 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 123914 592954
rect 123294 592634 123914 592718
rect 123294 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 123914 592634
rect 123294 556954 123914 592398
rect 123294 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 123914 556954
rect 123294 556634 123914 556718
rect 123294 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 123914 556634
rect 123294 520954 123914 556398
rect 123294 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 123914 520954
rect 123294 520634 123914 520718
rect 123294 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 123914 520634
rect 123294 484954 123914 520398
rect 123294 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 123914 484954
rect 123294 484634 123914 484718
rect 123294 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 123914 484634
rect 123294 448954 123914 484398
rect 123294 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 123914 448954
rect 123294 448634 123914 448718
rect 123294 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 123914 448634
rect 123294 412954 123914 448398
rect 123294 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 123914 412954
rect 123294 412634 123914 412718
rect 123294 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 123914 412634
rect 123294 376954 123914 412398
rect 123294 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 123914 376954
rect 123294 376634 123914 376718
rect 123294 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 123914 376634
rect 123294 340954 123914 376398
rect 123294 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 123914 340954
rect 123294 340634 123914 340718
rect 123294 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 123914 340634
rect 123294 304954 123914 340398
rect 123294 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 123914 304954
rect 123294 304634 123914 304718
rect 123294 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 123914 304634
rect 123294 268954 123914 304398
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 196954 123914 232398
rect 123294 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 123914 196954
rect 123294 196634 123914 196718
rect 123294 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 123914 196634
rect 123294 160954 123914 196398
rect 123294 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 123914 160954
rect 123294 160634 123914 160718
rect 123294 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 123914 160634
rect 123294 142000 123914 160398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 142000 128414 164898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 637954 132914 673398
rect 132294 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 132914 637954
rect 132294 637634 132914 637718
rect 132294 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 132914 637634
rect 132294 601954 132914 637398
rect 132294 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 132914 601954
rect 132294 601634 132914 601718
rect 132294 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 132914 601634
rect 132294 565954 132914 601398
rect 132294 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 132914 565954
rect 132294 565634 132914 565718
rect 132294 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 132914 565634
rect 132294 529954 132914 565398
rect 132294 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 132914 529954
rect 132294 529634 132914 529718
rect 132294 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 132914 529634
rect 132294 493954 132914 529398
rect 132294 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 132914 493954
rect 132294 493634 132914 493718
rect 132294 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 132914 493634
rect 132294 457954 132914 493398
rect 132294 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 132914 457954
rect 132294 457634 132914 457718
rect 132294 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 132914 457634
rect 132294 421954 132914 457398
rect 132294 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 132914 421954
rect 132294 421634 132914 421718
rect 132294 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 132914 421634
rect 132294 385954 132914 421398
rect 132294 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 132914 385954
rect 132294 385634 132914 385718
rect 132294 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 132914 385634
rect 132294 349954 132914 385398
rect 132294 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 132914 349954
rect 132294 349634 132914 349718
rect 132294 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 132914 349634
rect 132294 313954 132914 349398
rect 132294 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 132914 313954
rect 132294 313634 132914 313718
rect 132294 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 132914 313634
rect 132294 277954 132914 313398
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 205954 132914 241398
rect 132294 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 132914 205954
rect 132294 205634 132914 205718
rect 132294 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 132914 205634
rect 132294 169954 132914 205398
rect 132294 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 132914 169954
rect 132294 169634 132914 169718
rect 132294 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 132914 169634
rect 132294 142000 132914 169398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 642454 137414 677898
rect 136794 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 137414 642454
rect 136794 642134 137414 642218
rect 136794 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 137414 642134
rect 136794 606454 137414 641898
rect 136794 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 137414 606454
rect 136794 606134 137414 606218
rect 136794 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 137414 606134
rect 136794 570454 137414 605898
rect 136794 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 137414 570454
rect 136794 570134 137414 570218
rect 136794 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 137414 570134
rect 136794 534454 137414 569898
rect 136794 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 137414 534454
rect 136794 534134 137414 534218
rect 136794 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 137414 534134
rect 136794 498454 137414 533898
rect 136794 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 137414 498454
rect 136794 498134 137414 498218
rect 136794 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 137414 498134
rect 136794 462454 137414 497898
rect 136794 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 137414 462454
rect 136794 462134 137414 462218
rect 136794 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 137414 462134
rect 136794 426454 137414 461898
rect 136794 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 137414 426454
rect 136794 426134 137414 426218
rect 136794 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 137414 426134
rect 136794 390454 137414 425898
rect 136794 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 137414 390454
rect 136794 390134 137414 390218
rect 136794 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 137414 390134
rect 136794 354454 137414 389898
rect 136794 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 137414 354454
rect 136794 354134 137414 354218
rect 136794 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 137414 354134
rect 136794 318454 137414 353898
rect 136794 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 137414 318454
rect 136794 318134 137414 318218
rect 136794 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 137414 318134
rect 136794 282454 137414 317898
rect 136794 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 137414 282454
rect 136794 282134 137414 282218
rect 136794 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 137414 282134
rect 136794 246454 137414 281898
rect 136794 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 137414 246454
rect 136794 246134 137414 246218
rect 136794 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 137414 246134
rect 136794 210454 137414 245898
rect 136794 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 137414 210454
rect 136794 210134 137414 210218
rect 136794 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 137414 210134
rect 136794 174454 137414 209898
rect 136794 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 137414 174454
rect 136794 174134 137414 174218
rect 136794 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 137414 174134
rect 136794 142000 137414 173898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 646954 141914 682398
rect 141294 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 141914 646954
rect 141294 646634 141914 646718
rect 141294 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 141914 646634
rect 141294 610954 141914 646398
rect 141294 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 141914 610954
rect 141294 610634 141914 610718
rect 141294 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 141914 610634
rect 141294 574954 141914 610398
rect 141294 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 141914 574954
rect 141294 574634 141914 574718
rect 141294 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 141914 574634
rect 141294 538954 141914 574398
rect 141294 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 141914 538954
rect 141294 538634 141914 538718
rect 141294 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 141914 538634
rect 141294 502954 141914 538398
rect 141294 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 141914 502954
rect 141294 502634 141914 502718
rect 141294 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 141914 502634
rect 141294 466954 141914 502398
rect 141294 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 141914 466954
rect 141294 466634 141914 466718
rect 141294 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 141914 466634
rect 141294 430954 141914 466398
rect 141294 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 141914 430954
rect 141294 430634 141914 430718
rect 141294 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 141914 430634
rect 141294 394954 141914 430398
rect 141294 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 141914 394954
rect 141294 394634 141914 394718
rect 141294 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 141914 394634
rect 141294 358954 141914 394398
rect 141294 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 141914 358954
rect 141294 358634 141914 358718
rect 141294 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 141914 358634
rect 141294 322954 141914 358398
rect 141294 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 141914 322954
rect 141294 322634 141914 322718
rect 141294 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 141914 322634
rect 141294 286954 141914 322398
rect 141294 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 141914 286954
rect 141294 286634 141914 286718
rect 141294 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 141914 286634
rect 141294 250954 141914 286398
rect 141294 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 141914 250954
rect 141294 250634 141914 250718
rect 141294 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 141914 250634
rect 141294 214954 141914 250398
rect 141294 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 141914 214954
rect 141294 214634 141914 214718
rect 141294 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 141914 214634
rect 141294 178954 141914 214398
rect 141294 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 141914 178954
rect 141294 178634 141914 178718
rect 141294 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 141914 178634
rect 141294 142954 141914 178398
rect 141294 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 141914 142954
rect 141294 142634 141914 142718
rect 141294 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 141914 142634
rect 141294 142000 141914 142398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 142000 146414 146898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 655954 150914 691398
rect 150294 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 150914 655954
rect 150294 655634 150914 655718
rect 150294 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 150914 655634
rect 150294 619954 150914 655398
rect 150294 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 150914 619954
rect 150294 619634 150914 619718
rect 150294 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 150914 619634
rect 150294 583954 150914 619398
rect 150294 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 150914 583954
rect 150294 583634 150914 583718
rect 150294 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 150914 583634
rect 150294 547954 150914 583398
rect 150294 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 150914 547954
rect 150294 547634 150914 547718
rect 150294 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 150914 547634
rect 150294 511954 150914 547398
rect 150294 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 150914 511954
rect 150294 511634 150914 511718
rect 150294 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 150914 511634
rect 150294 475954 150914 511398
rect 150294 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 150914 475954
rect 150294 475634 150914 475718
rect 150294 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 150914 475634
rect 150294 439954 150914 475398
rect 150294 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 150914 439954
rect 150294 439634 150914 439718
rect 150294 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 150914 439634
rect 150294 403954 150914 439398
rect 150294 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 150914 403954
rect 150294 403634 150914 403718
rect 150294 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 150914 403634
rect 150294 367954 150914 403398
rect 150294 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 150914 367954
rect 150294 367634 150914 367718
rect 150294 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 150914 367634
rect 150294 331954 150914 367398
rect 150294 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 150914 331954
rect 150294 331634 150914 331718
rect 150294 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 150914 331634
rect 150294 295954 150914 331398
rect 150294 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 150914 295954
rect 150294 295634 150914 295718
rect 150294 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 150914 295634
rect 150294 259954 150914 295398
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 187954 150914 223398
rect 150294 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 150914 187954
rect 150294 187634 150914 187718
rect 150294 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 150914 187634
rect 150294 151954 150914 187398
rect 150294 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 150914 151954
rect 150294 151634 150914 151718
rect 150294 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 150914 151634
rect 150294 142000 150914 151398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 660454 155414 695898
rect 154794 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 155414 660454
rect 154794 660134 155414 660218
rect 154794 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 155414 660134
rect 154794 624454 155414 659898
rect 154794 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 155414 624454
rect 154794 624134 155414 624218
rect 154794 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 155414 624134
rect 154794 588454 155414 623898
rect 154794 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 155414 588454
rect 154794 588134 155414 588218
rect 154794 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 155414 588134
rect 154794 552454 155414 587898
rect 154794 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 155414 552454
rect 154794 552134 155414 552218
rect 154794 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 155414 552134
rect 154794 516454 155414 551898
rect 154794 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 155414 516454
rect 154794 516134 155414 516218
rect 154794 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 155414 516134
rect 154794 480454 155414 515898
rect 154794 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 155414 480454
rect 154794 480134 155414 480218
rect 154794 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 155414 480134
rect 154794 444454 155414 479898
rect 154794 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 155414 444454
rect 154794 444134 155414 444218
rect 154794 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 155414 444134
rect 154794 408454 155414 443898
rect 154794 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 155414 408454
rect 154794 408134 155414 408218
rect 154794 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 155414 408134
rect 154794 372454 155414 407898
rect 154794 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 155414 372454
rect 154794 372134 155414 372218
rect 154794 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 155414 372134
rect 154794 336454 155414 371898
rect 154794 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 155414 336454
rect 154794 336134 155414 336218
rect 154794 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 155414 336134
rect 154794 300454 155414 335898
rect 154794 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 155414 300454
rect 154794 300134 155414 300218
rect 154794 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 155414 300134
rect 154794 264454 155414 299898
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 192454 155414 227898
rect 154794 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 155414 192454
rect 154794 192134 155414 192218
rect 154794 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 155414 192134
rect 154794 156454 155414 191898
rect 154794 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 155414 156454
rect 154794 156134 155414 156218
rect 154794 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 155414 156134
rect 154794 142000 155414 155898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 628954 159914 664398
rect 159294 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 159914 628954
rect 159294 628634 159914 628718
rect 159294 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 159914 628634
rect 159294 592954 159914 628398
rect 159294 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 159914 592954
rect 159294 592634 159914 592718
rect 159294 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 159914 592634
rect 159294 556954 159914 592398
rect 159294 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 159914 556954
rect 159294 556634 159914 556718
rect 159294 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 159914 556634
rect 159294 520954 159914 556398
rect 159294 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 159914 520954
rect 159294 520634 159914 520718
rect 159294 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 159914 520634
rect 159294 484954 159914 520398
rect 159294 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 159914 484954
rect 159294 484634 159914 484718
rect 159294 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 159914 484634
rect 159294 448954 159914 484398
rect 159294 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 159914 448954
rect 159294 448634 159914 448718
rect 159294 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 159914 448634
rect 159294 412954 159914 448398
rect 159294 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 159914 412954
rect 159294 412634 159914 412718
rect 159294 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 159914 412634
rect 159294 376954 159914 412398
rect 159294 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 159914 376954
rect 159294 376634 159914 376718
rect 159294 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 159914 376634
rect 159294 340954 159914 376398
rect 159294 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 159914 340954
rect 159294 340634 159914 340718
rect 159294 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 159914 340634
rect 159294 304954 159914 340398
rect 159294 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 159914 304954
rect 159294 304634 159914 304718
rect 159294 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 159914 304634
rect 159294 268954 159914 304398
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 196954 159914 232398
rect 159294 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 159914 196954
rect 159294 196634 159914 196718
rect 159294 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 159914 196634
rect 159294 160954 159914 196398
rect 159294 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 159914 160954
rect 159294 160634 159914 160718
rect 159294 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 159914 160634
rect 159294 142000 159914 160398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 142000 164414 164898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 637954 168914 673398
rect 168294 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 168914 637954
rect 168294 637634 168914 637718
rect 168294 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 168914 637634
rect 168294 601954 168914 637398
rect 168294 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 168914 601954
rect 168294 601634 168914 601718
rect 168294 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 168914 601634
rect 168294 565954 168914 601398
rect 168294 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 168914 565954
rect 168294 565634 168914 565718
rect 168294 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 168914 565634
rect 168294 529954 168914 565398
rect 168294 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 168914 529954
rect 168294 529634 168914 529718
rect 168294 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 168914 529634
rect 168294 493954 168914 529398
rect 168294 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 168914 493954
rect 168294 493634 168914 493718
rect 168294 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 168914 493634
rect 168294 457954 168914 493398
rect 168294 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 168914 457954
rect 168294 457634 168914 457718
rect 168294 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 168914 457634
rect 168294 421954 168914 457398
rect 168294 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 168914 421954
rect 168294 421634 168914 421718
rect 168294 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 168914 421634
rect 168294 385954 168914 421398
rect 168294 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 168914 385954
rect 168294 385634 168914 385718
rect 168294 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 168914 385634
rect 168294 349954 168914 385398
rect 168294 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 168914 349954
rect 168294 349634 168914 349718
rect 168294 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 168914 349634
rect 168294 313954 168914 349398
rect 168294 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 168914 313954
rect 168294 313634 168914 313718
rect 168294 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 168914 313634
rect 168294 277954 168914 313398
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 205954 168914 241398
rect 168294 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 168914 205954
rect 168294 205634 168914 205718
rect 168294 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 168914 205634
rect 168294 169954 168914 205398
rect 168294 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 168914 169954
rect 168294 169634 168914 169718
rect 168294 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 168914 169634
rect 168294 142000 168914 169398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 642454 173414 677898
rect 172794 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 173414 642454
rect 172794 642134 173414 642218
rect 172794 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 173414 642134
rect 172794 606454 173414 641898
rect 172794 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 173414 606454
rect 172794 606134 173414 606218
rect 172794 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 173414 606134
rect 172794 570454 173414 605898
rect 172794 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 173414 570454
rect 172794 570134 173414 570218
rect 172794 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 173414 570134
rect 172794 534454 173414 569898
rect 172794 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 173414 534454
rect 172794 534134 173414 534218
rect 172794 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 173414 534134
rect 172794 498454 173414 533898
rect 172794 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 173414 498454
rect 172794 498134 173414 498218
rect 172794 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 173414 498134
rect 172794 462454 173414 497898
rect 172794 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 173414 462454
rect 172794 462134 173414 462218
rect 172794 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 173414 462134
rect 172794 426454 173414 461898
rect 172794 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 173414 426454
rect 172794 426134 173414 426218
rect 172794 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 173414 426134
rect 172794 390454 173414 425898
rect 172794 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 173414 390454
rect 172794 390134 173414 390218
rect 172794 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 173414 390134
rect 172794 354454 173414 389898
rect 172794 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 173414 354454
rect 172794 354134 173414 354218
rect 172794 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 173414 354134
rect 172794 318454 173414 353898
rect 172794 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 173414 318454
rect 172794 318134 173414 318218
rect 172794 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 173414 318134
rect 172794 282454 173414 317898
rect 172794 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 173414 282454
rect 172794 282134 173414 282218
rect 172794 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 173414 282134
rect 172794 246454 173414 281898
rect 172794 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 173414 246454
rect 172794 246134 173414 246218
rect 172794 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 173414 246134
rect 172794 210454 173414 245898
rect 172794 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 173414 210454
rect 172794 210134 173414 210218
rect 172794 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 173414 210134
rect 172794 174454 173414 209898
rect 172794 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 173414 174454
rect 172794 174134 173414 174218
rect 172794 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 173414 174134
rect 172794 142000 173414 173898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 646954 177914 682398
rect 177294 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 177914 646954
rect 177294 646634 177914 646718
rect 177294 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 177914 646634
rect 177294 610954 177914 646398
rect 177294 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 177914 610954
rect 177294 610634 177914 610718
rect 177294 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 177914 610634
rect 177294 574954 177914 610398
rect 177294 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 177914 574954
rect 177294 574634 177914 574718
rect 177294 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 177914 574634
rect 177294 538954 177914 574398
rect 177294 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 177914 538954
rect 177294 538634 177914 538718
rect 177294 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 177914 538634
rect 177294 502954 177914 538398
rect 177294 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 177914 502954
rect 177294 502634 177914 502718
rect 177294 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 177914 502634
rect 177294 466954 177914 502398
rect 177294 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 177914 466954
rect 177294 466634 177914 466718
rect 177294 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 177914 466634
rect 177294 430954 177914 466398
rect 177294 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 177914 430954
rect 177294 430634 177914 430718
rect 177294 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 177914 430634
rect 177294 394954 177914 430398
rect 177294 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 177914 394954
rect 177294 394634 177914 394718
rect 177294 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 177914 394634
rect 177294 358954 177914 394398
rect 177294 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 177914 358954
rect 177294 358634 177914 358718
rect 177294 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 177914 358634
rect 177294 322954 177914 358398
rect 177294 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 177914 322954
rect 177294 322634 177914 322718
rect 177294 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 177914 322634
rect 177294 286954 177914 322398
rect 177294 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 177914 286954
rect 177294 286634 177914 286718
rect 177294 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 177914 286634
rect 177294 250954 177914 286398
rect 177294 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 177914 250954
rect 177294 250634 177914 250718
rect 177294 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 177914 250634
rect 177294 214954 177914 250398
rect 177294 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 177914 214954
rect 177294 214634 177914 214718
rect 177294 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 177914 214634
rect 177294 178954 177914 214398
rect 177294 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 177914 178954
rect 177294 178634 177914 178718
rect 177294 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 177914 178634
rect 177294 142954 177914 178398
rect 177294 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 177914 142954
rect 177294 142634 177914 142718
rect 177294 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 177914 142634
rect 177294 142000 177914 142398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 655954 186914 691398
rect 186294 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 186914 655954
rect 186294 655634 186914 655718
rect 186294 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 186914 655634
rect 186294 619954 186914 655398
rect 186294 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 186914 619954
rect 186294 619634 186914 619718
rect 186294 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 186914 619634
rect 186294 583954 186914 619398
rect 186294 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 186914 583954
rect 186294 583634 186914 583718
rect 186294 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 186914 583634
rect 186294 547954 186914 583398
rect 186294 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 186914 547954
rect 186294 547634 186914 547718
rect 186294 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 186914 547634
rect 186294 511954 186914 547398
rect 186294 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 186914 511954
rect 186294 511634 186914 511718
rect 186294 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 186914 511634
rect 186294 475954 186914 511398
rect 186294 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 186914 475954
rect 186294 475634 186914 475718
rect 186294 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 186914 475634
rect 186294 439954 186914 475398
rect 186294 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 186914 439954
rect 186294 439634 186914 439718
rect 186294 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 186914 439634
rect 186294 403954 186914 439398
rect 186294 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 186914 403954
rect 186294 403634 186914 403718
rect 186294 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 186914 403634
rect 186294 367954 186914 403398
rect 186294 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 186914 367954
rect 186294 367634 186914 367718
rect 186294 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 186914 367634
rect 186294 331954 186914 367398
rect 186294 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 186914 331954
rect 186294 331634 186914 331718
rect 186294 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 186914 331634
rect 186294 295954 186914 331398
rect 186294 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 186914 295954
rect 186294 295634 186914 295718
rect 186294 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 186914 295634
rect 186294 259954 186914 295398
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 187954 186914 223398
rect 186294 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 186914 187954
rect 186294 187634 186914 187718
rect 186294 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 186914 187634
rect 186294 151954 186914 187398
rect 186294 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 186914 151954
rect 186294 151634 186914 151718
rect 186294 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 186914 151634
rect 186294 142000 186914 151398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 660454 191414 695898
rect 190794 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 191414 660454
rect 190794 660134 191414 660218
rect 190794 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 191414 660134
rect 190794 624454 191414 659898
rect 190794 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 191414 624454
rect 190794 624134 191414 624218
rect 190794 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 191414 624134
rect 190794 588454 191414 623898
rect 190794 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 191414 588454
rect 190794 588134 191414 588218
rect 190794 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 191414 588134
rect 190794 552454 191414 587898
rect 190794 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 191414 552454
rect 190794 552134 191414 552218
rect 190794 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 191414 552134
rect 190794 516454 191414 551898
rect 190794 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 191414 516454
rect 190794 516134 191414 516218
rect 190794 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 191414 516134
rect 190794 480454 191414 515898
rect 190794 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 191414 480454
rect 190794 480134 191414 480218
rect 190794 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 191414 480134
rect 190794 444454 191414 479898
rect 190794 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 191414 444454
rect 190794 444134 191414 444218
rect 190794 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 191414 444134
rect 190794 408454 191414 443898
rect 190794 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 191414 408454
rect 190794 408134 191414 408218
rect 190794 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 191414 408134
rect 190794 372454 191414 407898
rect 190794 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 191414 372454
rect 190794 372134 191414 372218
rect 190794 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 191414 372134
rect 190794 336454 191414 371898
rect 190794 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 191414 336454
rect 190794 336134 191414 336218
rect 190794 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 191414 336134
rect 190794 300454 191414 335898
rect 190794 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 191414 300454
rect 190794 300134 191414 300218
rect 190794 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 191414 300134
rect 190794 264454 191414 299898
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 192454 191414 227898
rect 190794 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 191414 192454
rect 190794 192134 191414 192218
rect 190794 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 191414 192134
rect 190794 156454 191414 191898
rect 190794 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 191414 156454
rect 190794 156134 191414 156218
rect 190794 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 191414 156134
rect 190794 142000 191414 155898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 628954 195914 664398
rect 195294 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 195914 628954
rect 195294 628634 195914 628718
rect 195294 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 195914 628634
rect 195294 592954 195914 628398
rect 195294 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 195914 592954
rect 195294 592634 195914 592718
rect 195294 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 195914 592634
rect 195294 556954 195914 592398
rect 195294 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 195914 556954
rect 195294 556634 195914 556718
rect 195294 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 195914 556634
rect 195294 520954 195914 556398
rect 195294 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 195914 520954
rect 195294 520634 195914 520718
rect 195294 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 195914 520634
rect 195294 484954 195914 520398
rect 195294 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 195914 484954
rect 195294 484634 195914 484718
rect 195294 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 195914 484634
rect 195294 448954 195914 484398
rect 195294 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 195914 448954
rect 195294 448634 195914 448718
rect 195294 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 195914 448634
rect 195294 412954 195914 448398
rect 195294 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 195914 412954
rect 195294 412634 195914 412718
rect 195294 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 195914 412634
rect 195294 376954 195914 412398
rect 195294 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 195914 376954
rect 195294 376634 195914 376718
rect 195294 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 195914 376634
rect 195294 340954 195914 376398
rect 195294 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 195914 340954
rect 195294 340634 195914 340718
rect 195294 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 195914 340634
rect 195294 304954 195914 340398
rect 195294 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 195914 304954
rect 195294 304634 195914 304718
rect 195294 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 195914 304634
rect 195294 268954 195914 304398
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 196954 195914 232398
rect 195294 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 195914 196954
rect 195294 196634 195914 196718
rect 195294 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 195914 196634
rect 195294 160954 195914 196398
rect 195294 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 195914 160954
rect 195294 160634 195914 160718
rect 195294 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 195914 160634
rect 195294 124954 195914 160398
rect 195294 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 195914 124954
rect 195294 124634 195914 124718
rect 195294 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 195914 124634
rect 114294 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 114914 115954
rect 114294 115634 114914 115718
rect 114294 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 114914 115634
rect 114294 79954 114914 115398
rect 139568 115954 139888 115986
rect 139568 115718 139610 115954
rect 139846 115718 139888 115954
rect 139568 115634 139888 115718
rect 139568 115398 139610 115634
rect 139846 115398 139888 115634
rect 139568 115366 139888 115398
rect 170288 115954 170608 115986
rect 170288 115718 170330 115954
rect 170566 115718 170608 115954
rect 170288 115634 170608 115718
rect 170288 115398 170330 115634
rect 170566 115398 170608 115634
rect 170288 115366 170608 115398
rect 124208 111454 124528 111486
rect 124208 111218 124250 111454
rect 124486 111218 124528 111454
rect 124208 111134 124528 111218
rect 124208 110898 124250 111134
rect 124486 110898 124528 111134
rect 124208 110866 124528 110898
rect 154928 111454 155248 111486
rect 154928 111218 154970 111454
rect 155206 111218 155248 111454
rect 154928 111134 155248 111218
rect 154928 110898 154970 111134
rect 155206 110898 155248 111134
rect 154928 110866 155248 110898
rect 185648 111454 185968 111486
rect 185648 111218 185690 111454
rect 185926 111218 185968 111454
rect 185648 111134 185968 111218
rect 185648 110898 185690 111134
rect 185926 110898 185968 111134
rect 185648 110866 185968 110898
rect 195294 88954 195914 124398
rect 195294 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 195914 88954
rect 195294 88634 195914 88718
rect 195294 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 195914 88634
rect 164371 80476 164437 80477
rect 164371 80412 164372 80476
rect 164436 80412 164437 80476
rect 164371 80411 164437 80412
rect 140819 80204 140885 80205
rect 140819 80140 140820 80204
rect 140884 80140 140885 80204
rect 140819 80139 140885 80140
rect 148363 80204 148429 80205
rect 148363 80140 148364 80204
rect 148428 80140 148429 80204
rect 148363 80139 148429 80140
rect 151307 80204 151373 80205
rect 151307 80140 151308 80204
rect 151372 80140 151373 80204
rect 151307 80139 151373 80140
rect 134195 80068 134261 80069
rect 134195 80066 134196 80068
rect 114294 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 114914 79954
rect 134014 80006 134196 80066
rect 131251 79932 131317 79933
rect 131251 79868 131252 79932
rect 131316 79868 131317 79932
rect 131251 79867 131317 79868
rect 131987 79932 132053 79933
rect 131987 79868 131988 79932
rect 132052 79868 132053 79932
rect 131987 79867 132053 79868
rect 132355 79932 132421 79933
rect 132355 79868 132356 79932
rect 132420 79868 132421 79932
rect 132355 79867 132421 79868
rect 132907 79932 132973 79933
rect 132907 79868 132908 79932
rect 132972 79868 132973 79932
rect 132907 79867 132973 79868
rect 114294 79634 114914 79718
rect 114294 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 114914 79634
rect 114294 43954 114914 79398
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 78000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 78000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 78000
rect 131067 73268 131133 73269
rect 131067 73204 131068 73268
rect 131132 73204 131133 73268
rect 131067 73203 131133 73204
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 131070 6493 131130 73203
rect 131254 35189 131314 79867
rect 131990 77893 132050 79867
rect 132358 78165 132418 79867
rect 132910 78165 132970 79867
rect 133091 79796 133157 79797
rect 133091 79732 133092 79796
rect 133156 79732 133157 79796
rect 133091 79731 133157 79732
rect 132355 78164 132421 78165
rect 132355 78100 132356 78164
rect 132420 78100 132421 78164
rect 132355 78099 132421 78100
rect 132907 78164 132973 78165
rect 132907 78100 132908 78164
rect 132972 78100 132973 78164
rect 132907 78099 132973 78100
rect 131987 77892 132053 77893
rect 131987 77828 131988 77892
rect 132052 77828 132053 77892
rect 131987 77827 132053 77828
rect 131619 77212 131685 77213
rect 131619 77148 131620 77212
rect 131684 77148 131685 77212
rect 131619 77147 131685 77148
rect 131622 72453 131682 77147
rect 131619 72452 131685 72453
rect 131619 72388 131620 72452
rect 131684 72388 131685 72452
rect 131619 72387 131685 72388
rect 132294 61954 132914 78000
rect 132294 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 132914 61954
rect 132294 61634 132914 61718
rect 132294 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 132914 61634
rect 131251 35188 131317 35189
rect 131251 35124 131252 35188
rect 131316 35124 131317 35188
rect 131251 35123 131317 35124
rect 132294 25954 132914 61398
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 131067 6492 131133 6493
rect 131067 6428 131068 6492
rect 131132 6428 131133 6492
rect 131067 6427 131133 6428
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 -5146 132914 25398
rect 133094 6357 133154 79731
rect 133275 75852 133341 75853
rect 133275 75788 133276 75852
rect 133340 75788 133341 75852
rect 133275 75787 133341 75788
rect 133091 6356 133157 6357
rect 133091 6292 133092 6356
rect 133156 6292 133157 6356
rect 133091 6291 133157 6292
rect 133278 6221 133338 75787
rect 134014 7717 134074 80006
rect 134195 80004 134196 80006
rect 134260 80004 134261 80068
rect 134195 80003 134261 80004
rect 134379 79932 134445 79933
rect 134379 79868 134380 79932
rect 134444 79868 134445 79932
rect 134379 79867 134445 79868
rect 135299 79932 135365 79933
rect 135299 79868 135300 79932
rect 135364 79868 135365 79932
rect 135299 79867 135365 79868
rect 136219 79932 136285 79933
rect 136219 79868 136220 79932
rect 136284 79868 136285 79932
rect 136219 79867 136285 79868
rect 137691 79932 137757 79933
rect 137691 79868 137692 79932
rect 137756 79868 137757 79932
rect 137691 79867 137757 79868
rect 137875 79932 137941 79933
rect 137875 79868 137876 79932
rect 137940 79868 137941 79932
rect 137875 79867 137941 79868
rect 138979 79932 139045 79933
rect 138979 79868 138980 79932
rect 139044 79868 139045 79932
rect 138979 79867 139045 79868
rect 139347 79932 139413 79933
rect 139347 79868 139348 79932
rect 139412 79868 139413 79932
rect 139347 79867 139413 79868
rect 134195 79796 134261 79797
rect 134195 79732 134196 79796
rect 134260 79732 134261 79796
rect 134195 79731 134261 79732
rect 134198 8941 134258 79731
rect 134195 8940 134261 8941
rect 134195 8876 134196 8940
rect 134260 8876 134261 8940
rect 134195 8875 134261 8876
rect 134011 7716 134077 7717
rect 134011 7652 134012 7716
rect 134076 7652 134077 7716
rect 134011 7651 134077 7652
rect 134382 7581 134442 79867
rect 134931 79796 134997 79797
rect 134931 79732 134932 79796
rect 134996 79732 134997 79796
rect 134931 79731 134997 79732
rect 134934 78709 134994 79731
rect 134931 78708 134997 78709
rect 134931 78644 134932 78708
rect 134996 78644 134997 78708
rect 134931 78643 134997 78644
rect 135302 7853 135362 79867
rect 135483 79796 135549 79797
rect 135483 79732 135484 79796
rect 135548 79794 135549 79796
rect 135851 79796 135917 79797
rect 135548 79734 135730 79794
rect 135548 79732 135549 79734
rect 135483 79731 135549 79732
rect 135483 77348 135549 77349
rect 135483 77284 135484 77348
rect 135548 77284 135549 77348
rect 135483 77283 135549 77284
rect 135486 7989 135546 77283
rect 135670 22677 135730 79734
rect 135851 79732 135852 79796
rect 135916 79732 135917 79796
rect 135851 79731 135917 79732
rect 135854 73813 135914 79731
rect 136222 78709 136282 79867
rect 136587 78844 136653 78845
rect 136587 78780 136588 78844
rect 136652 78780 136653 78844
rect 136587 78779 136653 78780
rect 136219 78708 136285 78709
rect 136219 78644 136220 78708
rect 136284 78644 136285 78708
rect 136219 78643 136285 78644
rect 136590 75445 136650 78779
rect 137694 78709 137754 79867
rect 137507 78708 137573 78709
rect 137507 78644 137508 78708
rect 137572 78644 137573 78708
rect 137507 78643 137573 78644
rect 137691 78708 137757 78709
rect 137691 78644 137692 78708
rect 137756 78644 137757 78708
rect 137691 78643 137757 78644
rect 136587 75444 136653 75445
rect 136587 75380 136588 75444
rect 136652 75380 136653 75444
rect 136587 75379 136653 75380
rect 135851 73812 135917 73813
rect 135851 73748 135852 73812
rect 135916 73748 135917 73812
rect 135851 73747 135917 73748
rect 136794 66454 137414 78000
rect 136794 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 137414 66454
rect 136794 66134 137414 66218
rect 136794 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 137414 66134
rect 136794 30454 137414 65898
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 135667 22676 135733 22677
rect 135667 22612 135668 22676
rect 135732 22612 135733 22676
rect 135667 22611 135733 22612
rect 135483 7988 135549 7989
rect 135483 7924 135484 7988
rect 135548 7924 135549 7988
rect 135483 7923 135549 7924
rect 135299 7852 135365 7853
rect 135299 7788 135300 7852
rect 135364 7788 135365 7852
rect 135299 7787 135365 7788
rect 134379 7580 134445 7581
rect 134379 7516 134380 7580
rect 134444 7516 134445 7580
rect 134379 7515 134445 7516
rect 133275 6220 133341 6221
rect 133275 6156 133276 6220
rect 133340 6156 133341 6220
rect 133275 6155 133341 6156
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 -6106 137414 29898
rect 137510 10301 137570 78643
rect 137878 77893 137938 79867
rect 138427 79796 138493 79797
rect 138427 79732 138428 79796
rect 138492 79732 138493 79796
rect 138427 79731 138493 79732
rect 138059 78844 138125 78845
rect 138059 78780 138060 78844
rect 138124 78780 138125 78844
rect 138059 78779 138125 78780
rect 137875 77892 137941 77893
rect 137875 77828 137876 77892
rect 137940 77828 137941 77892
rect 137875 77827 137941 77828
rect 137507 10300 137573 10301
rect 137507 10236 137508 10300
rect 137572 10236 137573 10300
rect 137507 10235 137573 10236
rect 138062 3365 138122 78779
rect 138243 78708 138309 78709
rect 138243 78644 138244 78708
rect 138308 78644 138309 78708
rect 138243 78643 138309 78644
rect 138246 10437 138306 78643
rect 138430 72725 138490 79731
rect 138982 78981 139042 79867
rect 138979 78980 139045 78981
rect 138979 78916 138980 78980
rect 139044 78916 139045 78980
rect 138979 78915 139045 78916
rect 139163 78164 139229 78165
rect 139163 78100 139164 78164
rect 139228 78100 139229 78164
rect 139163 78099 139229 78100
rect 138427 72724 138493 72725
rect 138427 72660 138428 72724
rect 138492 72660 138493 72724
rect 138427 72659 138493 72660
rect 139166 20365 139226 78099
rect 139350 76533 139410 79867
rect 139715 79796 139781 79797
rect 139715 79732 139716 79796
rect 139780 79732 139781 79796
rect 139715 79731 139781 79732
rect 139531 78708 139597 78709
rect 139531 78644 139532 78708
rect 139596 78644 139597 78708
rect 139531 78643 139597 78644
rect 139347 76532 139413 76533
rect 139347 76468 139348 76532
rect 139412 76468 139413 76532
rect 139347 76467 139413 76468
rect 139163 20364 139229 20365
rect 139163 20300 139164 20364
rect 139228 20300 139229 20364
rect 139163 20299 139229 20300
rect 139534 11661 139594 78643
rect 139531 11660 139597 11661
rect 139531 11596 139532 11660
rect 139596 11596 139597 11660
rect 139531 11595 139597 11596
rect 138243 10436 138309 10437
rect 138243 10372 138244 10436
rect 138308 10372 138309 10436
rect 138243 10371 138309 10372
rect 139718 9077 139778 79731
rect 140635 77348 140701 77349
rect 140635 77284 140636 77348
rect 140700 77284 140701 77348
rect 140635 77283 140701 77284
rect 140638 23085 140698 77283
rect 140635 23084 140701 23085
rect 140635 23020 140636 23084
rect 140700 23020 140701 23084
rect 140635 23019 140701 23020
rect 139715 9076 139781 9077
rect 139715 9012 139716 9076
rect 139780 9012 139781 9076
rect 139715 9011 139781 9012
rect 140822 3365 140882 80139
rect 143211 80068 143277 80069
rect 143211 80004 143212 80068
rect 143276 80004 143277 80068
rect 143211 80003 143277 80004
rect 141371 79932 141437 79933
rect 141371 79868 141372 79932
rect 141436 79868 141437 79932
rect 141371 79867 141437 79868
rect 142659 79932 142725 79933
rect 142659 79868 142660 79932
rect 142724 79868 142725 79932
rect 142659 79867 142725 79868
rect 141003 79796 141069 79797
rect 141003 79732 141004 79796
rect 141068 79732 141069 79796
rect 141003 79731 141069 79732
rect 141006 77621 141066 79731
rect 141374 78709 141434 79867
rect 141371 78708 141437 78709
rect 141371 78644 141372 78708
rect 141436 78644 141437 78708
rect 141371 78643 141437 78644
rect 141003 77620 141069 77621
rect 141003 77556 141004 77620
rect 141068 77556 141069 77620
rect 141003 77555 141069 77556
rect 141003 76668 141069 76669
rect 141003 76604 141004 76668
rect 141068 76604 141069 76668
rect 141003 76603 141069 76604
rect 141006 3637 141066 76603
rect 141294 70954 141914 78000
rect 142662 76669 142722 79867
rect 142843 77484 142909 77485
rect 142843 77420 142844 77484
rect 142908 77420 142909 77484
rect 142843 77419 142909 77420
rect 142659 76668 142725 76669
rect 142659 76604 142660 76668
rect 142724 76604 142725 76668
rect 142659 76603 142725 76604
rect 141294 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 141914 70954
rect 141294 70634 141914 70718
rect 141294 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 141914 70634
rect 141294 34954 141914 70398
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141003 3636 141069 3637
rect 141003 3572 141004 3636
rect 141068 3572 141069 3636
rect 141003 3571 141069 3572
rect 138059 3364 138125 3365
rect 138059 3300 138060 3364
rect 138124 3300 138125 3364
rect 138059 3299 138125 3300
rect 140819 3364 140885 3365
rect 140819 3300 140820 3364
rect 140884 3300 140885 3364
rect 140819 3299 140885 3300
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 -7066 141914 34398
rect 142846 18733 142906 77419
rect 143027 77348 143093 77349
rect 143027 77284 143028 77348
rect 143092 77284 143093 77348
rect 143027 77283 143093 77284
rect 142843 18732 142909 18733
rect 142843 18668 142844 18732
rect 142908 18668 142909 18732
rect 142843 18667 142909 18668
rect 143030 4997 143090 77283
rect 143027 4996 143093 4997
rect 143027 4932 143028 4996
rect 143092 4932 143093 4996
rect 143027 4931 143093 4932
rect 143214 4861 143274 80003
rect 143947 79932 144013 79933
rect 143947 79868 143948 79932
rect 144012 79868 144013 79932
rect 143947 79867 144013 79868
rect 144683 79932 144749 79933
rect 144683 79868 144684 79932
rect 144748 79868 144749 79932
rect 144683 79867 144749 79868
rect 145235 79932 145301 79933
rect 145235 79868 145236 79932
rect 145300 79868 145301 79932
rect 145235 79867 145301 79868
rect 146891 79932 146957 79933
rect 146891 79868 146892 79932
rect 146956 79868 146957 79932
rect 146891 79867 146957 79868
rect 148179 79932 148245 79933
rect 148179 79868 148180 79932
rect 148244 79868 148245 79932
rect 148179 79867 148245 79868
rect 143395 79796 143461 79797
rect 143395 79732 143396 79796
rect 143460 79732 143461 79796
rect 143395 79731 143461 79732
rect 143211 4860 143277 4861
rect 143211 4796 143212 4860
rect 143276 4796 143277 4860
rect 143211 4795 143277 4796
rect 143398 3501 143458 79731
rect 143950 76669 144010 79867
rect 144131 79796 144197 79797
rect 144131 79732 144132 79796
rect 144196 79732 144197 79796
rect 144131 79731 144197 79732
rect 143947 76668 144013 76669
rect 143947 76604 143948 76668
rect 144012 76604 144013 76668
rect 143947 76603 144013 76604
rect 144134 57221 144194 79731
rect 144499 77620 144565 77621
rect 144499 77556 144500 77620
rect 144564 77556 144565 77620
rect 144499 77555 144565 77556
rect 144315 77484 144381 77485
rect 144315 77420 144316 77484
rect 144380 77420 144381 77484
rect 144315 77419 144381 77420
rect 144318 68509 144378 77419
rect 144315 68508 144381 68509
rect 144315 68444 144316 68508
rect 144380 68444 144381 68508
rect 144315 68443 144381 68444
rect 144502 66877 144562 77555
rect 144686 75853 144746 79867
rect 145238 77485 145298 79867
rect 146523 79796 146589 79797
rect 146523 79732 146524 79796
rect 146588 79732 146589 79796
rect 146523 79731 146589 79732
rect 145235 77484 145301 77485
rect 145235 77420 145236 77484
rect 145300 77420 145301 77484
rect 145235 77419 145301 77420
rect 145419 77484 145485 77485
rect 145419 77420 145420 77484
rect 145484 77420 145485 77484
rect 145419 77419 145485 77420
rect 145235 77348 145301 77349
rect 145235 77284 145236 77348
rect 145300 77284 145301 77348
rect 145235 77283 145301 77284
rect 144683 75852 144749 75853
rect 144683 75788 144684 75852
rect 144748 75788 144749 75852
rect 144683 75787 144749 75788
rect 144499 66876 144565 66877
rect 144499 66812 144500 66876
rect 144564 66812 144565 66876
rect 144499 66811 144565 66812
rect 145238 63069 145298 77283
rect 145235 63068 145301 63069
rect 145235 63004 145236 63068
rect 145300 63004 145301 63068
rect 145235 63003 145301 63004
rect 144131 57220 144197 57221
rect 144131 57156 144132 57220
rect 144196 57156 144197 57220
rect 144131 57155 144197 57156
rect 145422 25533 145482 77419
rect 145603 76804 145669 76805
rect 145603 76740 145604 76804
rect 145668 76740 145669 76804
rect 145603 76739 145669 76740
rect 145419 25532 145485 25533
rect 145419 25468 145420 25532
rect 145484 25468 145485 25532
rect 145419 25467 145485 25468
rect 145606 20501 145666 76739
rect 145794 75454 146414 78000
rect 146526 76669 146586 79731
rect 146894 77349 146954 79867
rect 147075 79796 147141 79797
rect 147075 79732 147076 79796
rect 147140 79732 147141 79796
rect 147075 79731 147141 79732
rect 146891 77348 146957 77349
rect 146891 77284 146892 77348
rect 146956 77284 146957 77348
rect 146891 77283 146957 77284
rect 146523 76668 146589 76669
rect 146523 76604 146524 76668
rect 146588 76604 146589 76668
rect 146523 76603 146589 76604
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145603 20500 145669 20501
rect 145603 20436 145604 20500
rect 145668 20436 145669 20500
rect 145603 20435 145669 20436
rect 143395 3500 143461 3501
rect 143395 3436 143396 3500
rect 143460 3436 143461 3500
rect 143395 3435 143461 3436
rect 145794 3454 146414 38898
rect 147078 34237 147138 79731
rect 147443 77484 147509 77485
rect 147443 77420 147444 77484
rect 147508 77420 147509 77484
rect 147443 77419 147509 77420
rect 147259 77348 147325 77349
rect 147259 77284 147260 77348
rect 147324 77284 147325 77348
rect 147259 77283 147325 77284
rect 147075 34236 147141 34237
rect 147075 34172 147076 34236
rect 147140 34172 147141 34236
rect 147075 34171 147141 34172
rect 147262 23357 147322 77283
rect 147259 23356 147325 23357
rect 147259 23292 147260 23356
rect 147324 23292 147325 23356
rect 147259 23291 147325 23292
rect 147446 6085 147506 77419
rect 148182 76669 148242 79867
rect 148179 76668 148245 76669
rect 148179 76604 148180 76668
rect 148244 76604 148245 76668
rect 148179 76603 148245 76604
rect 148366 18597 148426 80139
rect 149099 79932 149165 79933
rect 149099 79868 149100 79932
rect 149164 79868 149165 79932
rect 149099 79867 149165 79868
rect 149467 79932 149533 79933
rect 149467 79868 149468 79932
rect 149532 79868 149533 79932
rect 149467 79867 149533 79868
rect 150755 79932 150821 79933
rect 150755 79868 150756 79932
rect 150820 79868 150821 79932
rect 150755 79867 150821 79868
rect 151123 79932 151189 79933
rect 151123 79868 151124 79932
rect 151188 79868 151189 79932
rect 151123 79867 151189 79868
rect 148731 79796 148797 79797
rect 148731 79732 148732 79796
rect 148796 79732 148797 79796
rect 148731 79731 148797 79732
rect 148547 75988 148613 75989
rect 148547 75924 148548 75988
rect 148612 75924 148613 75988
rect 148547 75923 148613 75924
rect 148363 18596 148429 18597
rect 148363 18532 148364 18596
rect 148428 18532 148429 18596
rect 148363 18531 148429 18532
rect 148550 10437 148610 75923
rect 148547 10436 148613 10437
rect 148547 10372 148548 10436
rect 148612 10372 148613 10436
rect 148547 10371 148613 10372
rect 147443 6084 147509 6085
rect 147443 6020 147444 6084
rect 147508 6020 147509 6084
rect 147443 6019 147509 6020
rect 148734 4045 148794 79731
rect 148915 76124 148981 76125
rect 148915 76060 148916 76124
rect 148980 76060 148981 76124
rect 148915 76059 148981 76060
rect 148731 4044 148797 4045
rect 148731 3980 148732 4044
rect 148796 3980 148797 4044
rect 148731 3979 148797 3980
rect 148918 3909 148978 76059
rect 149102 75989 149162 79867
rect 149470 76125 149530 79867
rect 149835 79796 149901 79797
rect 149835 79732 149836 79796
rect 149900 79732 149901 79796
rect 149835 79731 149901 79732
rect 149651 76668 149717 76669
rect 149651 76604 149652 76668
rect 149716 76604 149717 76668
rect 149651 76603 149717 76604
rect 149467 76124 149533 76125
rect 149467 76060 149468 76124
rect 149532 76060 149533 76124
rect 149467 76059 149533 76060
rect 149099 75988 149165 75989
rect 149099 75924 149100 75988
rect 149164 75924 149165 75988
rect 149099 75923 149165 75924
rect 149654 12069 149714 76603
rect 149651 12068 149717 12069
rect 149651 12004 149652 12068
rect 149716 12004 149717 12068
rect 149651 12003 149717 12004
rect 149838 6765 149898 79731
rect 150758 78301 150818 79867
rect 150755 78300 150821 78301
rect 150755 78236 150756 78300
rect 150820 78236 150821 78300
rect 150755 78235 150821 78236
rect 150019 75988 150085 75989
rect 150019 75924 150020 75988
rect 150084 75924 150085 75988
rect 150019 75923 150085 75924
rect 150022 6901 150082 75923
rect 150294 43954 150914 78000
rect 151126 75989 151186 79867
rect 151123 75988 151189 75989
rect 151123 75924 151124 75988
rect 151188 75924 151189 75988
rect 151123 75923 151189 75924
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 151310 28525 151370 80139
rect 163819 80068 163885 80069
rect 163819 80004 163820 80068
rect 163884 80004 163885 80068
rect 163819 80003 163885 80004
rect 151675 79932 151741 79933
rect 151675 79868 151676 79932
rect 151740 79868 151741 79932
rect 151675 79867 151741 79868
rect 152227 79932 152293 79933
rect 152227 79868 152228 79932
rect 152292 79868 152293 79932
rect 152963 79932 153029 79933
rect 152963 79930 152964 79932
rect 152227 79867 152293 79868
rect 152598 79870 152964 79930
rect 151491 75988 151557 75989
rect 151491 75924 151492 75988
rect 151556 75924 151557 75988
rect 151491 75923 151557 75924
rect 151307 28524 151373 28525
rect 151307 28460 151308 28524
rect 151372 28460 151373 28524
rect 151307 28459 151373 28460
rect 151494 11933 151554 75923
rect 151491 11932 151557 11933
rect 151491 11868 151492 11932
rect 151556 11868 151557 11932
rect 151491 11867 151557 11868
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150019 6900 150085 6901
rect 150019 6836 150020 6900
rect 150084 6836 150085 6900
rect 150019 6835 150085 6836
rect 149835 6764 149901 6765
rect 149835 6700 149836 6764
rect 149900 6700 149901 6764
rect 149835 6699 149901 6700
rect 148915 3908 148981 3909
rect 148915 3844 148916 3908
rect 148980 3844 148981 3908
rect 148915 3843 148981 3844
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 -1306 150914 7398
rect 151678 6629 151738 79867
rect 152230 75989 152290 79867
rect 152411 79796 152477 79797
rect 152411 79732 152412 79796
rect 152476 79732 152477 79796
rect 152411 79731 152477 79732
rect 152227 75988 152293 75989
rect 152227 75924 152228 75988
rect 152292 75924 152293 75988
rect 152227 75923 152293 75924
rect 152414 23221 152474 79731
rect 152411 23220 152477 23221
rect 152411 23156 152412 23220
rect 152476 23156 152477 23220
rect 152411 23155 152477 23156
rect 152598 14517 152658 79870
rect 152963 79868 152964 79870
rect 153028 79868 153029 79932
rect 152963 79867 153029 79868
rect 153699 79932 153765 79933
rect 153699 79868 153700 79932
rect 153764 79868 153765 79932
rect 153699 79867 153765 79868
rect 154067 79932 154133 79933
rect 154067 79868 154068 79932
rect 154132 79868 154133 79932
rect 154067 79867 154133 79868
rect 154619 79932 154685 79933
rect 154619 79868 154620 79932
rect 154684 79868 154685 79932
rect 154619 79867 154685 79868
rect 155539 79932 155605 79933
rect 155539 79868 155540 79932
rect 155604 79868 155605 79932
rect 155539 79867 155605 79868
rect 155907 79932 155973 79933
rect 155907 79868 155908 79932
rect 155972 79868 155973 79932
rect 155907 79867 155973 79868
rect 156459 79932 156525 79933
rect 156459 79868 156460 79932
rect 156524 79868 156525 79932
rect 156459 79867 156525 79868
rect 157011 79932 157077 79933
rect 157011 79868 157012 79932
rect 157076 79868 157077 79932
rect 157011 79867 157077 79868
rect 157931 79932 157997 79933
rect 157931 79868 157932 79932
rect 157996 79868 157997 79932
rect 157931 79867 157997 79868
rect 158299 79932 158365 79933
rect 158299 79868 158300 79932
rect 158364 79868 158365 79932
rect 158299 79867 158365 79868
rect 160507 79932 160573 79933
rect 160507 79868 160508 79932
rect 160572 79868 160573 79932
rect 161243 79932 161309 79933
rect 161243 79930 161244 79932
rect 160507 79867 160573 79868
rect 161062 79870 161244 79930
rect 152779 76124 152845 76125
rect 152779 76060 152780 76124
rect 152844 76060 152845 76124
rect 152779 76059 152845 76060
rect 152595 14516 152661 14517
rect 152595 14452 152596 14516
rect 152660 14452 152661 14516
rect 152595 14451 152661 14452
rect 151675 6628 151741 6629
rect 151675 6564 151676 6628
rect 151740 6564 151741 6628
rect 151675 6563 151741 6564
rect 152782 6357 152842 76059
rect 153702 75989 153762 79867
rect 153883 77076 153949 77077
rect 153883 77012 153884 77076
rect 153948 77012 153949 77076
rect 153883 77011 153949 77012
rect 152963 75988 153029 75989
rect 152963 75924 152964 75988
rect 153028 75924 153029 75988
rect 152963 75923 153029 75924
rect 153699 75988 153765 75989
rect 153699 75924 153700 75988
rect 153764 75924 153765 75988
rect 153699 75923 153765 75924
rect 152966 6493 153026 75923
rect 153886 9213 153946 77011
rect 153883 9212 153949 9213
rect 153883 9148 153884 9212
rect 153948 9148 153949 9212
rect 153883 9147 153949 9148
rect 154070 9077 154130 79867
rect 154622 75989 154682 79867
rect 155542 79117 155602 79867
rect 155539 79116 155605 79117
rect 155539 79052 155540 79116
rect 155604 79052 155605 79116
rect 155539 79051 155605 79052
rect 154251 75988 154317 75989
rect 154251 75924 154252 75988
rect 154316 75924 154317 75988
rect 154251 75923 154317 75924
rect 154619 75988 154685 75989
rect 154619 75924 154620 75988
rect 154684 75924 154685 75988
rect 154619 75923 154685 75924
rect 154067 9076 154133 9077
rect 154067 9012 154068 9076
rect 154132 9012 154133 9076
rect 154067 9011 154133 9012
rect 154254 8941 154314 75923
rect 154794 48454 155414 78000
rect 155910 75037 155970 79867
rect 155907 75036 155973 75037
rect 155907 74972 155908 75036
rect 155972 74972 155973 75036
rect 155907 74971 155973 74972
rect 156462 73813 156522 79867
rect 156643 79796 156709 79797
rect 156643 79732 156644 79796
rect 156708 79732 156709 79796
rect 156643 79731 156709 79732
rect 156827 79796 156893 79797
rect 156827 79732 156828 79796
rect 156892 79732 156893 79796
rect 156827 79731 156893 79732
rect 156646 78981 156706 79731
rect 156643 78980 156709 78981
rect 156643 78916 156644 78980
rect 156708 78916 156709 78980
rect 156643 78915 156709 78916
rect 156830 76261 156890 79731
rect 156827 76260 156893 76261
rect 156827 76196 156828 76260
rect 156892 76196 156893 76260
rect 156827 76195 156893 76196
rect 156643 76124 156709 76125
rect 156643 76060 156644 76124
rect 156708 76060 156709 76124
rect 156643 76059 156709 76060
rect 156459 73812 156525 73813
rect 156459 73748 156460 73812
rect 156524 73748 156525 73812
rect 156459 73747 156525 73748
rect 156646 71637 156706 76059
rect 157014 74357 157074 79867
rect 157934 76941 157994 79867
rect 158115 79796 158181 79797
rect 158115 79732 158116 79796
rect 158180 79732 158181 79796
rect 158115 79731 158181 79732
rect 157931 76940 157997 76941
rect 157931 76876 157932 76940
rect 157996 76876 157997 76940
rect 157931 76875 157997 76876
rect 157011 74356 157077 74357
rect 157011 74292 157012 74356
rect 157076 74292 157077 74356
rect 157011 74291 157077 74292
rect 158118 71773 158178 79731
rect 158302 72589 158362 79867
rect 158483 79660 158549 79661
rect 158483 79596 158484 79660
rect 158548 79596 158549 79660
rect 158483 79595 158549 79596
rect 158299 72588 158365 72589
rect 158299 72524 158300 72588
rect 158364 72524 158365 72588
rect 158299 72523 158365 72524
rect 158115 71772 158181 71773
rect 158115 71708 158116 71772
rect 158180 71708 158181 71772
rect 158115 71707 158181 71708
rect 156643 71636 156709 71637
rect 156643 71572 156644 71636
rect 156708 71572 156709 71636
rect 156643 71571 156709 71572
rect 158486 68373 158546 79595
rect 158851 78980 158917 78981
rect 158851 78916 158852 78980
rect 158916 78916 158917 78980
rect 158851 78915 158917 78916
rect 158854 71501 158914 78915
rect 158851 71500 158917 71501
rect 158851 71436 158852 71500
rect 158916 71436 158917 71500
rect 158851 71435 158917 71436
rect 158483 68372 158549 68373
rect 158483 68308 158484 68372
rect 158548 68308 158549 68372
rect 158483 68307 158549 68308
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154251 8940 154317 8941
rect 154251 8876 154252 8940
rect 154316 8876 154317 8940
rect 154251 8875 154317 8876
rect 152963 6492 153029 6493
rect 152963 6428 152964 6492
rect 153028 6428 153029 6492
rect 152963 6427 153029 6428
rect 152779 6356 152845 6357
rect 152779 6292 152780 6356
rect 152844 6292 152845 6356
rect 152779 6291 152845 6292
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 52954 159914 78000
rect 160510 76941 160570 79867
rect 160691 78844 160757 78845
rect 160691 78780 160692 78844
rect 160756 78780 160757 78844
rect 160691 78779 160757 78780
rect 160507 76940 160573 76941
rect 160507 76876 160508 76940
rect 160572 76876 160573 76940
rect 160507 76875 160573 76876
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 160694 10301 160754 78779
rect 160875 78708 160941 78709
rect 160875 78644 160876 78708
rect 160940 78644 160941 78708
rect 160875 78643 160941 78644
rect 160878 74629 160938 78643
rect 160875 74628 160941 74629
rect 160875 74564 160876 74628
rect 160940 74564 160941 74628
rect 160875 74563 160941 74564
rect 161062 48925 161122 79870
rect 161243 79868 161244 79870
rect 161308 79868 161309 79932
rect 161243 79867 161309 79868
rect 161611 79932 161677 79933
rect 161611 79868 161612 79932
rect 161676 79868 161677 79932
rect 161611 79867 161677 79868
rect 161979 79932 162045 79933
rect 161979 79868 161980 79932
rect 162044 79868 162045 79932
rect 161979 79867 162045 79868
rect 162347 79932 162413 79933
rect 162347 79868 162348 79932
rect 162412 79868 162413 79932
rect 162347 79867 162413 79868
rect 162715 79932 162781 79933
rect 162715 79868 162716 79932
rect 162780 79868 162781 79932
rect 162715 79867 162781 79868
rect 163635 79932 163701 79933
rect 163635 79868 163636 79932
rect 163700 79868 163701 79932
rect 163635 79867 163701 79868
rect 161614 78709 161674 79867
rect 161982 78845 162042 79867
rect 162163 79116 162229 79117
rect 162163 79052 162164 79116
rect 162228 79052 162229 79116
rect 162163 79051 162229 79052
rect 161979 78844 162045 78845
rect 161979 78780 161980 78844
rect 162044 78780 162045 78844
rect 161979 78779 162045 78780
rect 161611 78708 161677 78709
rect 161611 78644 161612 78708
rect 161676 78644 161677 78708
rect 161611 78643 161677 78644
rect 161243 77348 161309 77349
rect 161243 77284 161244 77348
rect 161308 77284 161309 77348
rect 161243 77283 161309 77284
rect 161246 74221 161306 77283
rect 161427 74628 161493 74629
rect 161427 74564 161428 74628
rect 161492 74564 161493 74628
rect 161427 74563 161493 74564
rect 161243 74220 161309 74221
rect 161243 74156 161244 74220
rect 161308 74156 161309 74220
rect 161243 74155 161309 74156
rect 161430 71365 161490 74563
rect 161427 71364 161493 71365
rect 161427 71300 161428 71364
rect 161492 71300 161493 71364
rect 161427 71299 161493 71300
rect 161059 48924 161125 48925
rect 161059 48860 161060 48924
rect 161124 48860 161125 48924
rect 161059 48859 161125 48860
rect 162166 20093 162226 79051
rect 162350 78981 162410 79867
rect 162531 79660 162597 79661
rect 162531 79596 162532 79660
rect 162596 79596 162597 79660
rect 162531 79595 162597 79596
rect 162347 78980 162413 78981
rect 162347 78916 162348 78980
rect 162412 78916 162413 78980
rect 162347 78915 162413 78916
rect 162347 78708 162413 78709
rect 162347 78644 162348 78708
rect 162412 78644 162413 78708
rect 162347 78643 162413 78644
rect 162350 20229 162410 78643
rect 162347 20228 162413 20229
rect 162347 20164 162348 20228
rect 162412 20164 162413 20228
rect 162347 20163 162413 20164
rect 162163 20092 162229 20093
rect 162163 20028 162164 20092
rect 162228 20028 162229 20092
rect 162163 20027 162229 20028
rect 162534 11797 162594 79595
rect 162531 11796 162597 11797
rect 162531 11732 162532 11796
rect 162596 11732 162597 11796
rect 162531 11731 162597 11732
rect 162718 11661 162778 79867
rect 163083 79660 163149 79661
rect 163083 79596 163084 79660
rect 163148 79596 163149 79660
rect 163083 79595 163149 79596
rect 163086 78709 163146 79595
rect 163638 79117 163698 79867
rect 163635 79116 163701 79117
rect 163635 79052 163636 79116
rect 163700 79052 163701 79116
rect 163635 79051 163701 79052
rect 163267 78844 163333 78845
rect 163267 78780 163268 78844
rect 163332 78780 163333 78844
rect 163267 78779 163333 78780
rect 163083 78708 163149 78709
rect 163083 78644 163084 78708
rect 163148 78644 163149 78708
rect 163083 78643 163149 78644
rect 163270 33965 163330 78779
rect 163451 78708 163517 78709
rect 163451 78644 163452 78708
rect 163516 78644 163517 78708
rect 163822 78706 163882 80003
rect 164374 79933 164434 80411
rect 177987 80340 178053 80341
rect 177987 80276 177988 80340
rect 178052 80276 178053 80340
rect 177987 80275 178053 80276
rect 168603 80204 168669 80205
rect 168603 80140 168604 80204
rect 168668 80140 168669 80204
rect 168603 80139 168669 80140
rect 164371 79932 164437 79933
rect 164371 79868 164372 79932
rect 164436 79868 164437 79932
rect 164371 79867 164437 79868
rect 164923 79932 164989 79933
rect 164923 79868 164924 79932
rect 164988 79930 164989 79932
rect 166579 79932 166645 79933
rect 164988 79870 165354 79930
rect 164988 79868 164989 79870
rect 164923 79867 164989 79868
rect 164003 79796 164069 79797
rect 164003 79732 164004 79796
rect 164068 79732 164069 79796
rect 164003 79731 164069 79732
rect 164006 78981 164066 79731
rect 164923 79660 164989 79661
rect 164923 79596 164924 79660
rect 164988 79596 164989 79660
rect 164923 79595 164989 79596
rect 164003 78980 164069 78981
rect 164003 78916 164004 78980
rect 164068 78916 164069 78980
rect 164003 78915 164069 78916
rect 163451 78643 163517 78644
rect 163638 78646 163882 78706
rect 163454 34101 163514 78643
rect 163451 34100 163517 34101
rect 163451 34036 163452 34100
rect 163516 34036 163517 34100
rect 163451 34035 163517 34036
rect 163267 33964 163333 33965
rect 163267 33900 163268 33964
rect 163332 33900 163333 33964
rect 163267 33899 163333 33900
rect 163638 31381 163698 78646
rect 163794 57454 164414 78000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163635 31380 163701 31381
rect 163635 31316 163636 31380
rect 163700 31316 163701 31380
rect 163635 31315 163701 31316
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 162715 11660 162781 11661
rect 162715 11596 162716 11660
rect 162780 11596 162781 11660
rect 162715 11595 162781 11596
rect 160691 10300 160757 10301
rect 160691 10236 160692 10300
rect 160756 10236 160757 10300
rect 160691 10235 160757 10236
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 -4186 164414 20898
rect 164926 17509 164986 79595
rect 165107 78708 165173 78709
rect 165107 78644 165108 78708
rect 165172 78644 165173 78708
rect 165107 78643 165173 78644
rect 165110 17645 165170 78643
rect 165294 17781 165354 79870
rect 166579 79868 166580 79932
rect 166644 79868 166645 79932
rect 166579 79867 166645 79868
rect 166763 79932 166829 79933
rect 166763 79868 166764 79932
rect 166828 79868 166829 79932
rect 166763 79867 166829 79868
rect 167315 79932 167381 79933
rect 167315 79868 167316 79932
rect 167380 79868 167381 79932
rect 167315 79867 167381 79868
rect 168051 79932 168117 79933
rect 168051 79868 168052 79932
rect 168116 79868 168117 79932
rect 168051 79867 168117 79868
rect 166395 79660 166461 79661
rect 166395 79596 166396 79660
rect 166460 79596 166461 79660
rect 166395 79595 166461 79596
rect 165475 78708 165541 78709
rect 165475 78644 165476 78708
rect 165540 78644 165541 78708
rect 165475 78643 165541 78644
rect 165291 17780 165357 17781
rect 165291 17716 165292 17780
rect 165356 17716 165357 17780
rect 165291 17715 165357 17716
rect 165107 17644 165173 17645
rect 165107 17580 165108 17644
rect 165172 17580 165173 17644
rect 165107 17579 165173 17580
rect 164923 17508 164989 17509
rect 164923 17444 164924 17508
rect 164988 17444 164989 17508
rect 164923 17443 164989 17444
rect 165478 6221 165538 78643
rect 166211 78300 166277 78301
rect 166211 78236 166212 78300
rect 166276 78236 166277 78300
rect 166211 78235 166277 78236
rect 166214 31245 166274 78235
rect 166211 31244 166277 31245
rect 166211 31180 166212 31244
rect 166276 31180 166277 31244
rect 166211 31179 166277 31180
rect 166398 28389 166458 79595
rect 166582 78845 166642 79867
rect 166766 79661 166826 79867
rect 166763 79660 166829 79661
rect 166763 79596 166764 79660
rect 166828 79596 166829 79660
rect 166763 79595 166829 79596
rect 166579 78844 166645 78845
rect 166579 78780 166580 78844
rect 166644 78780 166645 78844
rect 166579 78779 166645 78780
rect 166763 78844 166829 78845
rect 166763 78780 166764 78844
rect 166828 78780 166829 78844
rect 166763 78779 166829 78780
rect 166579 78708 166645 78709
rect 166579 78644 166580 78708
rect 166644 78644 166645 78708
rect 166579 78643 166645 78644
rect 166395 28388 166461 28389
rect 166395 28324 166396 28388
rect 166460 28324 166461 28388
rect 166395 28323 166461 28324
rect 166582 17237 166642 78643
rect 166766 17373 166826 78779
rect 167318 78165 167378 79867
rect 167867 79660 167933 79661
rect 167867 79596 167868 79660
rect 167932 79596 167933 79660
rect 167867 79595 167933 79596
rect 167683 78980 167749 78981
rect 167683 78916 167684 78980
rect 167748 78916 167749 78980
rect 167683 78915 167749 78916
rect 167499 78708 167565 78709
rect 167499 78644 167500 78708
rect 167564 78644 167565 78708
rect 167499 78643 167565 78644
rect 167315 78164 167381 78165
rect 167315 78100 167316 78164
rect 167380 78100 167381 78164
rect 167315 78099 167381 78100
rect 167502 31109 167562 78643
rect 167686 69597 167746 78915
rect 167683 69596 167749 69597
rect 167683 69532 167684 69596
rect 167748 69532 167749 69596
rect 167683 69531 167749 69532
rect 167870 68237 167930 79595
rect 168054 72453 168114 79867
rect 168606 79525 168666 80139
rect 171363 80068 171429 80069
rect 171363 80004 171364 80068
rect 171428 80004 171429 80068
rect 171363 80003 171429 80004
rect 174307 80068 174373 80069
rect 174307 80004 174308 80068
rect 174372 80004 174373 80068
rect 177067 80068 177133 80069
rect 174307 80003 174373 80004
rect 175782 80006 176210 80066
rect 169155 79932 169221 79933
rect 169155 79868 169156 79932
rect 169220 79868 169221 79932
rect 169155 79867 169221 79868
rect 169523 79932 169589 79933
rect 169523 79868 169524 79932
rect 169588 79868 169589 79932
rect 169523 79867 169589 79868
rect 170075 79932 170141 79933
rect 170075 79868 170076 79932
rect 170140 79868 170141 79932
rect 170075 79867 170141 79868
rect 168603 79524 168669 79525
rect 168603 79460 168604 79524
rect 168668 79460 168669 79524
rect 168603 79459 168669 79460
rect 168051 72452 168117 72453
rect 168051 72388 168052 72452
rect 168116 72388 168117 72452
rect 168051 72387 168117 72388
rect 167867 68236 167933 68237
rect 167867 68172 167868 68236
rect 167932 68172 167933 68236
rect 167867 68171 167933 68172
rect 168294 61954 168914 78000
rect 169158 75989 169218 79867
rect 169155 75988 169221 75989
rect 169155 75924 169156 75988
rect 169220 75924 169221 75988
rect 169155 75923 169221 75924
rect 168294 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 168914 61954
rect 168294 61634 168914 61718
rect 168294 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 168914 61634
rect 167499 31108 167565 31109
rect 167499 31044 167500 31108
rect 167564 31044 167565 31108
rect 167499 31043 167565 31044
rect 168294 25954 168914 61398
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 166763 17372 166829 17373
rect 166763 17308 166764 17372
rect 166828 17308 166829 17372
rect 166763 17307 166829 17308
rect 166579 17236 166645 17237
rect 166579 17172 166580 17236
rect 166644 17172 166645 17236
rect 166579 17171 166645 17172
rect 165475 6220 165541 6221
rect 165475 6156 165476 6220
rect 165540 6156 165541 6220
rect 165475 6155 165541 6156
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 -5146 168914 25398
rect 169526 21317 169586 79867
rect 169707 78708 169773 78709
rect 169707 78644 169708 78708
rect 169772 78644 169773 78708
rect 169707 78643 169773 78644
rect 169710 71229 169770 78643
rect 170078 75989 170138 79867
rect 170627 79796 170693 79797
rect 170627 79732 170628 79796
rect 170692 79732 170693 79796
rect 170627 79731 170693 79732
rect 170443 79524 170509 79525
rect 170443 79460 170444 79524
rect 170508 79460 170509 79524
rect 170443 79459 170509 79460
rect 170259 77892 170325 77893
rect 170259 77828 170260 77892
rect 170324 77828 170325 77892
rect 170259 77827 170325 77828
rect 170075 75988 170141 75989
rect 170075 75924 170076 75988
rect 170140 75924 170141 75988
rect 170075 75923 170141 75924
rect 169707 71228 169773 71229
rect 169707 71164 169708 71228
rect 169772 71164 169773 71228
rect 169707 71163 169773 71164
rect 170262 22949 170322 77827
rect 170446 77213 170506 79459
rect 170443 77212 170509 77213
rect 170443 77148 170444 77212
rect 170508 77148 170509 77212
rect 170443 77147 170509 77148
rect 170630 71093 170690 79731
rect 170995 78708 171061 78709
rect 170995 78644 170996 78708
rect 171060 78644 171061 78708
rect 170995 78643 171061 78644
rect 170811 75988 170877 75989
rect 170811 75924 170812 75988
rect 170876 75924 170877 75988
rect 170811 75923 170877 75924
rect 170627 71092 170693 71093
rect 170627 71028 170628 71092
rect 170692 71028 170693 71092
rect 170627 71027 170693 71028
rect 170814 24309 170874 75923
rect 170811 24308 170877 24309
rect 170811 24244 170812 24308
rect 170876 24244 170877 24308
rect 170811 24243 170877 24244
rect 170259 22948 170325 22949
rect 170259 22884 170260 22948
rect 170324 22884 170325 22948
rect 170259 22883 170325 22884
rect 170998 22813 171058 78643
rect 171366 76125 171426 80003
rect 172099 79932 172165 79933
rect 172099 79868 172100 79932
rect 172164 79868 172165 79932
rect 172099 79867 172165 79868
rect 173387 79932 173453 79933
rect 173387 79868 173388 79932
rect 173452 79868 173453 79932
rect 173387 79867 173453 79868
rect 173755 79932 173821 79933
rect 173755 79868 173756 79932
rect 173820 79868 173821 79932
rect 173755 79867 173821 79868
rect 174123 79932 174189 79933
rect 174123 79868 174124 79932
rect 174188 79868 174189 79932
rect 174123 79867 174189 79868
rect 171547 79796 171613 79797
rect 171547 79732 171548 79796
rect 171612 79732 171613 79796
rect 171547 79731 171613 79732
rect 171363 76124 171429 76125
rect 171363 76060 171364 76124
rect 171428 76060 171429 76124
rect 171363 76059 171429 76060
rect 171550 75989 171610 79731
rect 171915 79524 171981 79525
rect 171915 79460 171916 79524
rect 171980 79460 171981 79524
rect 171915 79459 171981 79460
rect 171731 78708 171797 78709
rect 171731 78644 171732 78708
rect 171796 78644 171797 78708
rect 171731 78643 171797 78644
rect 171547 75988 171613 75989
rect 171547 75924 171548 75988
rect 171612 75924 171613 75988
rect 171547 75923 171613 75924
rect 170995 22812 171061 22813
rect 170995 22748 170996 22812
rect 171060 22748 171061 22812
rect 170995 22747 171061 22748
rect 169523 21316 169589 21317
rect 169523 21252 169524 21316
rect 169588 21252 169589 21316
rect 169523 21251 169589 21252
rect 171734 19957 171794 78643
rect 171918 61573 171978 79459
rect 172102 78573 172162 79867
rect 173390 79525 173450 79867
rect 173387 79524 173453 79525
rect 173387 79460 173388 79524
rect 173452 79460 173453 79524
rect 173387 79459 173453 79460
rect 172099 78572 172165 78573
rect 172099 78508 172100 78572
rect 172164 78508 172165 78572
rect 172099 78507 172165 78508
rect 172099 78436 172165 78437
rect 172099 78372 172100 78436
rect 172164 78372 172165 78436
rect 172099 78371 172165 78372
rect 171915 61572 171981 61573
rect 171915 61508 171916 61572
rect 171980 61508 171981 61572
rect 171915 61507 171981 61508
rect 172102 22677 172162 78371
rect 172794 66454 173414 78000
rect 173571 77348 173637 77349
rect 173571 77284 173572 77348
rect 173636 77284 173637 77348
rect 173571 77283 173637 77284
rect 172794 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 173414 66454
rect 172794 66134 173414 66218
rect 172794 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 173414 66134
rect 172794 30454 173414 65898
rect 173574 33829 173634 77283
rect 173571 33828 173637 33829
rect 173571 33764 173572 33828
rect 173636 33764 173637 33828
rect 173571 33763 173637 33764
rect 173758 30973 173818 79867
rect 174126 77893 174186 79867
rect 174310 78165 174370 80003
rect 175782 79933 175842 80006
rect 174675 79932 174741 79933
rect 174675 79868 174676 79932
rect 174740 79868 174741 79932
rect 174675 79867 174741 79868
rect 175227 79932 175293 79933
rect 175227 79868 175228 79932
rect 175292 79868 175293 79932
rect 175227 79867 175293 79868
rect 175779 79932 175845 79933
rect 175779 79868 175780 79932
rect 175844 79868 175845 79932
rect 175779 79867 175845 79868
rect 174491 79796 174557 79797
rect 174491 79732 174492 79796
rect 174556 79732 174557 79796
rect 174491 79731 174557 79732
rect 174307 78164 174373 78165
rect 174307 78100 174308 78164
rect 174372 78100 174373 78164
rect 174307 78099 174373 78100
rect 174123 77892 174189 77893
rect 174123 77828 174124 77892
rect 174188 77828 174189 77892
rect 174123 77827 174189 77828
rect 174494 73541 174554 79731
rect 174678 78437 174738 79867
rect 174859 79116 174925 79117
rect 174859 79052 174860 79116
rect 174924 79052 174925 79116
rect 174859 79051 174925 79052
rect 174675 78436 174741 78437
rect 174675 78372 174676 78436
rect 174740 78372 174741 78436
rect 174675 78371 174741 78372
rect 174675 78164 174741 78165
rect 174675 78100 174676 78164
rect 174740 78100 174741 78164
rect 174675 78099 174741 78100
rect 174491 73540 174557 73541
rect 174491 73476 174492 73540
rect 174556 73476 174557 73540
rect 174491 73475 174557 73476
rect 173755 30972 173821 30973
rect 173755 30908 173756 30972
rect 173820 30908 173821 30972
rect 173755 30907 173821 30908
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172099 22676 172165 22677
rect 172099 22612 172100 22676
rect 172164 22612 172165 22676
rect 172099 22611 172165 22612
rect 171731 19956 171797 19957
rect 171731 19892 171732 19956
rect 171796 19892 171797 19956
rect 171731 19891 171797 19892
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 -6106 173414 29898
rect 174678 24173 174738 78099
rect 174862 62933 174922 79051
rect 175230 78709 175290 79867
rect 175227 78708 175293 78709
rect 175227 78644 175228 78708
rect 175292 78644 175293 78708
rect 175227 78643 175293 78644
rect 175963 78708 176029 78709
rect 175963 78644 175964 78708
rect 176028 78644 176029 78708
rect 175963 78643 176029 78644
rect 175966 75989 176026 78643
rect 175963 75988 176029 75989
rect 175963 75924 175964 75988
rect 176028 75924 176029 75988
rect 175963 75923 176029 75924
rect 174859 62932 174925 62933
rect 174859 62868 174860 62932
rect 174924 62868 174925 62932
rect 174859 62867 174925 62868
rect 176150 62797 176210 80006
rect 177067 80004 177068 80068
rect 177132 80004 177133 80068
rect 177067 80003 177133 80004
rect 176331 79796 176397 79797
rect 176331 79732 176332 79796
rect 176396 79732 176397 79796
rect 176331 79731 176397 79732
rect 176147 62796 176213 62797
rect 176147 62732 176148 62796
rect 176212 62732 176213 62796
rect 176147 62731 176213 62732
rect 176334 61437 176394 79731
rect 176515 78436 176581 78437
rect 176515 78372 176516 78436
rect 176580 78372 176581 78436
rect 176515 78371 176581 78372
rect 176331 61436 176397 61437
rect 176331 61372 176332 61436
rect 176396 61372 176397 61436
rect 176331 61371 176397 61372
rect 176518 46205 176578 78371
rect 176883 77892 176949 77893
rect 176883 77828 176884 77892
rect 176948 77828 176949 77892
rect 176883 77827 176949 77828
rect 176515 46204 176581 46205
rect 176515 46140 176516 46204
rect 176580 46140 176581 46204
rect 176515 46139 176581 46140
rect 174675 24172 174741 24173
rect 174675 24108 174676 24172
rect 174740 24108 174741 24172
rect 174675 24107 174741 24108
rect 176886 3365 176946 77827
rect 177070 77621 177130 80003
rect 177990 79661 178050 80275
rect 178539 79932 178605 79933
rect 178539 79868 178540 79932
rect 178604 79868 178605 79932
rect 178539 79867 178605 79868
rect 177987 79660 178053 79661
rect 177987 79596 177988 79660
rect 178052 79596 178053 79660
rect 177987 79595 178053 79596
rect 178542 79253 178602 79867
rect 178539 79252 178605 79253
rect 178539 79188 178540 79252
rect 178604 79188 178605 79252
rect 178539 79187 178605 79188
rect 177067 77620 177133 77621
rect 177067 77556 177068 77620
rect 177132 77556 177133 77620
rect 177067 77555 177133 77556
rect 177067 76124 177133 76125
rect 177067 76060 177068 76124
rect 177132 76060 177133 76124
rect 177067 76059 177133 76060
rect 177070 3501 177130 76059
rect 177294 70954 177914 78000
rect 177294 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 177914 70954
rect 177294 70634 177914 70718
rect 177294 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 177914 70634
rect 177294 34954 177914 70398
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177067 3500 177133 3501
rect 177067 3436 177068 3500
rect 177132 3436 177133 3500
rect 177067 3435 177133 3436
rect 176883 3364 176949 3365
rect 176883 3300 176884 3364
rect 176948 3300 176949 3364
rect 176883 3299 176949 3300
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 75454 182414 78000
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 78000
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 78000
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 52954 195914 88398
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 637954 204914 673398
rect 204294 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 204914 637954
rect 204294 637634 204914 637718
rect 204294 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 204914 637634
rect 204294 601954 204914 637398
rect 204294 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 204914 601954
rect 204294 601634 204914 601718
rect 204294 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 204914 601634
rect 204294 565954 204914 601398
rect 204294 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 204914 565954
rect 204294 565634 204914 565718
rect 204294 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 204914 565634
rect 204294 529954 204914 565398
rect 204294 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 204914 529954
rect 204294 529634 204914 529718
rect 204294 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 204914 529634
rect 204294 493954 204914 529398
rect 204294 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 204914 493954
rect 204294 493634 204914 493718
rect 204294 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 204914 493634
rect 204294 457954 204914 493398
rect 204294 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 204914 457954
rect 204294 457634 204914 457718
rect 204294 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 204914 457634
rect 204294 421954 204914 457398
rect 204294 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 204914 421954
rect 204294 421634 204914 421718
rect 204294 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 204914 421634
rect 204294 385954 204914 421398
rect 204294 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 204914 385954
rect 204294 385634 204914 385718
rect 204294 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 204914 385634
rect 204294 349954 204914 385398
rect 204294 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 204914 349954
rect 204294 349634 204914 349718
rect 204294 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 204914 349634
rect 204294 313954 204914 349398
rect 204294 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 204914 313954
rect 204294 313634 204914 313718
rect 204294 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 204914 313634
rect 204294 277954 204914 313398
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 205954 204914 241398
rect 204294 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 204914 205954
rect 204294 205634 204914 205718
rect 204294 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 204914 205634
rect 204294 169954 204914 205398
rect 204294 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 204914 169954
rect 204294 169634 204914 169718
rect 204294 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 204914 169634
rect 204294 133954 204914 169398
rect 204294 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 204914 133954
rect 204294 133634 204914 133718
rect 204294 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 204914 133634
rect 204294 97954 204914 133398
rect 204294 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 204914 97954
rect 204294 97634 204914 97718
rect 204294 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 204914 97634
rect 204294 61954 204914 97398
rect 204294 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 204914 61954
rect 204294 61634 204914 61718
rect 204294 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 204914 61634
rect 204294 25954 204914 61398
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 642454 209414 677898
rect 208794 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 209414 642454
rect 208794 642134 209414 642218
rect 208794 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 209414 642134
rect 208794 606454 209414 641898
rect 208794 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 209414 606454
rect 208794 606134 209414 606218
rect 208794 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 209414 606134
rect 208794 570454 209414 605898
rect 208794 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 209414 570454
rect 208794 570134 209414 570218
rect 208794 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 209414 570134
rect 208794 534454 209414 569898
rect 208794 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 209414 534454
rect 208794 534134 209414 534218
rect 208794 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 209414 534134
rect 208794 498454 209414 533898
rect 208794 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 209414 498454
rect 208794 498134 209414 498218
rect 208794 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 209414 498134
rect 208794 462454 209414 497898
rect 208794 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 209414 462454
rect 208794 462134 209414 462218
rect 208794 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 209414 462134
rect 208794 426454 209414 461898
rect 208794 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 209414 426454
rect 208794 426134 209414 426218
rect 208794 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 209414 426134
rect 208794 390454 209414 425898
rect 208794 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 209414 390454
rect 208794 390134 209414 390218
rect 208794 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 209414 390134
rect 208794 354454 209414 389898
rect 208794 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 209414 354454
rect 208794 354134 209414 354218
rect 208794 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 209414 354134
rect 208794 318454 209414 353898
rect 208794 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 209414 318454
rect 208794 318134 209414 318218
rect 208794 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 209414 318134
rect 208794 282454 209414 317898
rect 208794 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 209414 282454
rect 208794 282134 209414 282218
rect 208794 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 209414 282134
rect 208794 246454 209414 281898
rect 208794 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 209414 246454
rect 208794 246134 209414 246218
rect 208794 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 209414 246134
rect 208794 210454 209414 245898
rect 208794 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 209414 210454
rect 208794 210134 209414 210218
rect 208794 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 209414 210134
rect 208794 174454 209414 209898
rect 208794 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 209414 174454
rect 208794 174134 209414 174218
rect 208794 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 209414 174134
rect 208794 138454 209414 173898
rect 208794 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 209414 138454
rect 208794 138134 209414 138218
rect 208794 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 209414 138134
rect 208794 102454 209414 137898
rect 208794 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 209414 102454
rect 208794 102134 209414 102218
rect 208794 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 209414 102134
rect 208794 66454 209414 101898
rect 208794 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 209414 66454
rect 208794 66134 209414 66218
rect 208794 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 209414 66134
rect 208794 30454 209414 65898
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 646954 213914 682398
rect 213294 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 213914 646954
rect 213294 646634 213914 646718
rect 213294 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 213914 646634
rect 213294 610954 213914 646398
rect 213294 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 213914 610954
rect 213294 610634 213914 610718
rect 213294 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 213914 610634
rect 213294 574954 213914 610398
rect 213294 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 213914 574954
rect 213294 574634 213914 574718
rect 213294 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 213914 574634
rect 213294 538954 213914 574398
rect 213294 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 213914 538954
rect 213294 538634 213914 538718
rect 213294 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 213914 538634
rect 213294 502954 213914 538398
rect 213294 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 213914 502954
rect 213294 502634 213914 502718
rect 213294 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 213914 502634
rect 213294 466954 213914 502398
rect 213294 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 213914 466954
rect 213294 466634 213914 466718
rect 213294 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 213914 466634
rect 213294 430954 213914 466398
rect 213294 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 213914 430954
rect 213294 430634 213914 430718
rect 213294 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 213914 430634
rect 213294 394954 213914 430398
rect 213294 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 213914 394954
rect 213294 394634 213914 394718
rect 213294 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 213914 394634
rect 213294 358954 213914 394398
rect 213294 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 213914 358954
rect 213294 358634 213914 358718
rect 213294 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 213914 358634
rect 213294 322954 213914 358398
rect 213294 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 213914 322954
rect 213294 322634 213914 322718
rect 213294 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 213914 322634
rect 213294 286954 213914 322398
rect 213294 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 213914 286954
rect 213294 286634 213914 286718
rect 213294 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 213914 286634
rect 213294 250954 213914 286398
rect 213294 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 213914 250954
rect 213294 250634 213914 250718
rect 213294 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 213914 250634
rect 213294 214954 213914 250398
rect 213294 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 213914 214954
rect 213294 214634 213914 214718
rect 213294 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 213914 214634
rect 213294 178954 213914 214398
rect 213294 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 213914 178954
rect 213294 178634 213914 178718
rect 213294 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 213914 178634
rect 213294 142954 213914 178398
rect 213294 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 213914 142954
rect 213294 142634 213914 142718
rect 213294 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 213914 142634
rect 213294 106954 213914 142398
rect 213294 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 213914 106954
rect 213294 106634 213914 106718
rect 213294 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 213914 106634
rect 213294 70954 213914 106398
rect 213294 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 213914 70954
rect 213294 70634 213914 70718
rect 213294 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 213914 70634
rect 213294 34954 213914 70398
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 655954 222914 691398
rect 222294 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 222914 655954
rect 222294 655634 222914 655718
rect 222294 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 222914 655634
rect 222294 619954 222914 655398
rect 222294 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 222914 619954
rect 222294 619634 222914 619718
rect 222294 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 222914 619634
rect 222294 583954 222914 619398
rect 222294 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 222914 583954
rect 222294 583634 222914 583718
rect 222294 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 222914 583634
rect 222294 547954 222914 583398
rect 222294 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 222914 547954
rect 222294 547634 222914 547718
rect 222294 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 222914 547634
rect 222294 511954 222914 547398
rect 222294 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 222914 511954
rect 222294 511634 222914 511718
rect 222294 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 222914 511634
rect 222294 475954 222914 511398
rect 222294 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 222914 475954
rect 222294 475634 222914 475718
rect 222294 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 222914 475634
rect 222294 439954 222914 475398
rect 222294 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 222914 439954
rect 222294 439634 222914 439718
rect 222294 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 222914 439634
rect 222294 403954 222914 439398
rect 222294 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 222914 403954
rect 222294 403634 222914 403718
rect 222294 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 222914 403634
rect 222294 367954 222914 403398
rect 222294 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 222914 367954
rect 222294 367634 222914 367718
rect 222294 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 222914 367634
rect 222294 331954 222914 367398
rect 222294 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 222914 331954
rect 222294 331634 222914 331718
rect 222294 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 222914 331634
rect 222294 295954 222914 331398
rect 222294 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 222914 295954
rect 222294 295634 222914 295718
rect 222294 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 222914 295634
rect 222294 259954 222914 295398
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 187954 222914 223398
rect 222294 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 222914 187954
rect 222294 187634 222914 187718
rect 222294 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 222914 187634
rect 222294 151954 222914 187398
rect 222294 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 222914 151954
rect 222294 151634 222914 151718
rect 222294 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 222914 151634
rect 222294 115954 222914 151398
rect 222294 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 222914 115954
rect 222294 115634 222914 115718
rect 222294 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 222914 115634
rect 222294 79954 222914 115398
rect 222294 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 222914 79954
rect 222294 79634 222914 79718
rect 222294 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 222914 79634
rect 222294 43954 222914 79398
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 660454 227414 695898
rect 226794 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 227414 660454
rect 226794 660134 227414 660218
rect 226794 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 227414 660134
rect 226794 624454 227414 659898
rect 226794 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 227414 624454
rect 226794 624134 227414 624218
rect 226794 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 227414 624134
rect 226794 588454 227414 623898
rect 226794 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 227414 588454
rect 226794 588134 227414 588218
rect 226794 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 227414 588134
rect 226794 552454 227414 587898
rect 226794 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 227414 552454
rect 226794 552134 227414 552218
rect 226794 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 227414 552134
rect 226794 516454 227414 551898
rect 226794 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 227414 516454
rect 226794 516134 227414 516218
rect 226794 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 227414 516134
rect 226794 480454 227414 515898
rect 226794 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 227414 480454
rect 226794 480134 227414 480218
rect 226794 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 227414 480134
rect 226794 444454 227414 479898
rect 226794 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 227414 444454
rect 226794 444134 227414 444218
rect 226794 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 227414 444134
rect 226794 408454 227414 443898
rect 226794 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 227414 408454
rect 226794 408134 227414 408218
rect 226794 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 227414 408134
rect 226794 372454 227414 407898
rect 226794 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 227414 372454
rect 226794 372134 227414 372218
rect 226794 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 227414 372134
rect 226794 336454 227414 371898
rect 226794 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 227414 336454
rect 226794 336134 227414 336218
rect 226794 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 227414 336134
rect 226794 300454 227414 335898
rect 226794 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 227414 300454
rect 226794 300134 227414 300218
rect 226794 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 227414 300134
rect 226794 264454 227414 299898
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 628954 231914 664398
rect 231294 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 231914 628954
rect 231294 628634 231914 628718
rect 231294 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 231914 628634
rect 231294 592954 231914 628398
rect 231294 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 231914 592954
rect 231294 592634 231914 592718
rect 231294 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 231914 592634
rect 231294 556954 231914 592398
rect 231294 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 231914 556954
rect 231294 556634 231914 556718
rect 231294 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 231914 556634
rect 231294 520954 231914 556398
rect 231294 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 231914 520954
rect 231294 520634 231914 520718
rect 231294 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 231914 520634
rect 231294 484954 231914 520398
rect 231294 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 231914 484954
rect 231294 484634 231914 484718
rect 231294 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 231914 484634
rect 231294 448954 231914 484398
rect 231294 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 231914 448954
rect 231294 448634 231914 448718
rect 231294 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 231914 448634
rect 231294 412954 231914 448398
rect 231294 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 231914 412954
rect 231294 412634 231914 412718
rect 231294 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 231914 412634
rect 231294 376954 231914 412398
rect 231294 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 231914 376954
rect 231294 376634 231914 376718
rect 231294 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 231914 376634
rect 231294 340954 231914 376398
rect 231294 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 231914 340954
rect 231294 340634 231914 340718
rect 231294 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 231914 340634
rect 231294 304954 231914 340398
rect 231294 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 231914 304954
rect 231294 304634 231914 304718
rect 231294 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 231914 304634
rect 231294 268954 231914 304398
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 637954 240914 673398
rect 240294 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 240914 637954
rect 240294 637634 240914 637718
rect 240294 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 240914 637634
rect 240294 601954 240914 637398
rect 240294 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 240914 601954
rect 240294 601634 240914 601718
rect 240294 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 240914 601634
rect 240294 565954 240914 601398
rect 240294 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 240914 565954
rect 240294 565634 240914 565718
rect 240294 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 240914 565634
rect 240294 529954 240914 565398
rect 240294 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 240914 529954
rect 240294 529634 240914 529718
rect 240294 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 240914 529634
rect 240294 493954 240914 529398
rect 240294 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 240914 493954
rect 240294 493634 240914 493718
rect 240294 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 240914 493634
rect 240294 457954 240914 493398
rect 240294 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 240914 457954
rect 240294 457634 240914 457718
rect 240294 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 240914 457634
rect 240294 421954 240914 457398
rect 240294 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 240914 421954
rect 240294 421634 240914 421718
rect 240294 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 240914 421634
rect 240294 385954 240914 421398
rect 240294 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 240914 385954
rect 240294 385634 240914 385718
rect 240294 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 240914 385634
rect 240294 349954 240914 385398
rect 240294 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 240914 349954
rect 240294 349634 240914 349718
rect 240294 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 240914 349634
rect 240294 313954 240914 349398
rect 240294 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 240914 313954
rect 240294 313634 240914 313718
rect 240294 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 240914 313634
rect 240294 277954 240914 313398
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 642454 245414 677898
rect 244794 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 245414 642454
rect 244794 642134 245414 642218
rect 244794 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 245414 642134
rect 244794 606454 245414 641898
rect 244794 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 245414 606454
rect 244794 606134 245414 606218
rect 244794 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 245414 606134
rect 244794 570454 245414 605898
rect 244794 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 245414 570454
rect 244794 570134 245414 570218
rect 244794 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 245414 570134
rect 244794 534454 245414 569898
rect 244794 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 245414 534454
rect 244794 534134 245414 534218
rect 244794 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 245414 534134
rect 244794 498454 245414 533898
rect 244794 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 245414 498454
rect 244794 498134 245414 498218
rect 244794 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 245414 498134
rect 244794 462454 245414 497898
rect 244794 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 245414 462454
rect 244794 462134 245414 462218
rect 244794 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 245414 462134
rect 244794 426454 245414 461898
rect 244794 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 245414 426454
rect 244794 426134 245414 426218
rect 244794 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 245414 426134
rect 244794 390454 245414 425898
rect 244794 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 245414 390454
rect 244794 390134 245414 390218
rect 244794 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 245414 390134
rect 244794 354454 245414 389898
rect 244794 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 245414 354454
rect 244794 354134 245414 354218
rect 244794 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 245414 354134
rect 244794 318454 245414 353898
rect 244794 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 245414 318454
rect 244794 318134 245414 318218
rect 244794 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 245414 318134
rect 244794 282454 245414 317898
rect 244794 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 245414 282454
rect 244794 282134 245414 282218
rect 244794 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 245414 282134
rect 244794 246454 245414 281898
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 646954 249914 682398
rect 249294 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 249914 646954
rect 249294 646634 249914 646718
rect 249294 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 249914 646634
rect 249294 610954 249914 646398
rect 249294 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 249914 610954
rect 249294 610634 249914 610718
rect 249294 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 249914 610634
rect 249294 574954 249914 610398
rect 249294 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 249914 574954
rect 249294 574634 249914 574718
rect 249294 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 249914 574634
rect 249294 538954 249914 574398
rect 249294 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 249914 538954
rect 249294 538634 249914 538718
rect 249294 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 249914 538634
rect 249294 502954 249914 538398
rect 249294 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 249914 502954
rect 249294 502634 249914 502718
rect 249294 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 249914 502634
rect 249294 466954 249914 502398
rect 249294 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 249914 466954
rect 249294 466634 249914 466718
rect 249294 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 249914 466634
rect 249294 430954 249914 466398
rect 249294 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 249914 430954
rect 249294 430634 249914 430718
rect 249294 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 249914 430634
rect 249294 394954 249914 430398
rect 249294 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 249914 394954
rect 249294 394634 249914 394718
rect 249294 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 249914 394634
rect 249294 358954 249914 394398
rect 249294 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 249914 358954
rect 249294 358634 249914 358718
rect 249294 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 249914 358634
rect 249294 322954 249914 358398
rect 249294 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 249914 322954
rect 249294 322634 249914 322718
rect 249294 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 249914 322634
rect 249294 286954 249914 322398
rect 249294 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 249914 286954
rect 249294 286634 249914 286718
rect 249294 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 249914 286634
rect 249294 250954 249914 286398
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 637954 276914 673398
rect 276294 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 276914 637954
rect 276294 637634 276914 637718
rect 276294 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 276914 637634
rect 276294 601954 276914 637398
rect 276294 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 276914 601954
rect 276294 601634 276914 601718
rect 276294 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 276914 601634
rect 276294 565954 276914 601398
rect 276294 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 276914 565954
rect 276294 565634 276914 565718
rect 276294 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 276914 565634
rect 276294 529954 276914 565398
rect 276294 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 276914 529954
rect 276294 529634 276914 529718
rect 276294 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 276914 529634
rect 276294 493954 276914 529398
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 280794 642454 281414 677898
rect 280794 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 281414 642454
rect 280794 642134 281414 642218
rect 280794 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 281414 642134
rect 280794 606454 281414 641898
rect 280794 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 281414 606454
rect 280794 606134 281414 606218
rect 280794 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 281414 606134
rect 280794 570454 281414 605898
rect 280794 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 281414 570454
rect 280794 570134 281414 570218
rect 280794 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 281414 570134
rect 280794 534454 281414 569898
rect 280794 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 281414 534454
rect 280794 534134 281414 534218
rect 280794 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 281414 534134
rect 280794 498454 281414 533898
rect 280794 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 281414 498454
rect 280794 498134 281414 498218
rect 280794 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 281414 498134
rect 280794 462454 281414 497898
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 285294 646954 285914 682398
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 610954 285914 646398
rect 285294 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 285914 610954
rect 285294 610634 285914 610718
rect 285294 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 285914 610634
rect 285294 574954 285914 610398
rect 285294 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 285914 574954
rect 285294 574634 285914 574718
rect 285294 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 285914 574634
rect 285294 538954 285914 574398
rect 285294 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 285914 538954
rect 285294 538634 285914 538718
rect 285294 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 285914 538634
rect 285294 502954 285914 538398
rect 285294 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 285914 502954
rect 285294 502634 285914 502718
rect 285294 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 285914 502634
rect 285294 466954 285914 502398
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 285294 250954 285914 286398
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 619954 294914 655398
rect 294294 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 294914 619954
rect 294294 619634 294914 619718
rect 294294 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 294914 619634
rect 294294 583954 294914 619398
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 511954 294914 547398
rect 294294 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 294914 511954
rect 294294 511634 294914 511718
rect 294294 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 294914 511634
rect 294294 475954 294914 511398
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 294294 259954 294914 295398
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 624454 299414 659898
rect 298794 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 299414 624454
rect 298794 624134 299414 624218
rect 298794 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 299414 624134
rect 298794 588454 299414 623898
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 298794 516454 299414 551898
rect 298794 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 299414 516454
rect 298794 516134 299414 516218
rect 298794 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 299414 516134
rect 298794 480454 299414 515898
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 298794 300454 299414 335898
rect 298794 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 299414 300454
rect 298794 300134 299414 300218
rect 298794 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 299414 300134
rect 298794 264454 299414 299898
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 192454 299414 227898
rect 298794 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 299414 192454
rect 298794 192134 299414 192218
rect 298794 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 299414 192134
rect 298794 156454 299414 191898
rect 298794 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 299414 156454
rect 298794 156134 299414 156218
rect 298794 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 299414 156134
rect 298794 120454 299414 155898
rect 298794 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 299414 120454
rect 298794 120134 299414 120218
rect 298794 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 299414 120134
rect 298794 84454 299414 119898
rect 298794 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 299414 84454
rect 298794 84134 299414 84218
rect 298794 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 299414 84134
rect 298794 48454 299414 83898
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298794 -2266 299414 11898
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 628954 303914 664398
rect 303294 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 303914 628954
rect 303294 628634 303914 628718
rect 303294 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 303914 628634
rect 303294 592954 303914 628398
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 520954 303914 556398
rect 303294 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 303914 520954
rect 303294 520634 303914 520718
rect 303294 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 303914 520634
rect 303294 484954 303914 520398
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 303294 304954 303914 340398
rect 303294 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 303914 304954
rect 303294 304634 303914 304718
rect 303294 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 303914 304634
rect 303294 268954 303914 304398
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 196954 303914 232398
rect 303294 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 303914 196954
rect 303294 196634 303914 196718
rect 303294 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 303914 196634
rect 303294 160954 303914 196398
rect 303294 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 303914 160954
rect 303294 160634 303914 160718
rect 303294 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 303914 160634
rect 303294 124954 303914 160398
rect 303294 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 303914 124954
rect 303294 124634 303914 124718
rect 303294 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 303914 124634
rect 303294 88954 303914 124398
rect 303294 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 303914 88954
rect 303294 88634 303914 88718
rect 303294 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 303914 88634
rect 303294 52954 303914 88398
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 312294 637954 312914 673398
rect 312294 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 312914 637954
rect 312294 637634 312914 637718
rect 312294 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 312914 637634
rect 312294 601954 312914 637398
rect 312294 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 312914 601954
rect 312294 601634 312914 601718
rect 312294 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 312914 601634
rect 312294 565954 312914 601398
rect 312294 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 312914 565954
rect 312294 565634 312914 565718
rect 312294 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 312914 565634
rect 312294 529954 312914 565398
rect 312294 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 312914 529954
rect 312294 529634 312914 529718
rect 312294 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 312914 529634
rect 312294 493954 312914 529398
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 313954 312914 349398
rect 312294 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 312914 313954
rect 312294 313634 312914 313718
rect 312294 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 312914 313634
rect 312294 277954 312914 313398
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 205954 312914 241398
rect 312294 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 312914 205954
rect 312294 205634 312914 205718
rect 312294 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 312914 205634
rect 312294 169954 312914 205398
rect 312294 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 312914 169954
rect 312294 169634 312914 169718
rect 312294 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 312914 169634
rect 312294 133954 312914 169398
rect 312294 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 312914 133954
rect 312294 133634 312914 133718
rect 312294 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 312914 133634
rect 312294 97954 312914 133398
rect 312294 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 312914 97954
rect 312294 97634 312914 97718
rect 312294 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 312914 97634
rect 312294 61954 312914 97398
rect 312294 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 312914 61954
rect 312294 61634 312914 61718
rect 312294 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 312914 61634
rect 312294 25954 312914 61398
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642454 317414 677898
rect 316794 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 317414 642454
rect 316794 642134 317414 642218
rect 316794 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 317414 642134
rect 316794 606454 317414 641898
rect 316794 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 317414 606454
rect 316794 606134 317414 606218
rect 316794 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 317414 606134
rect 316794 570454 317414 605898
rect 316794 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 317414 570454
rect 316794 570134 317414 570218
rect 316794 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 317414 570134
rect 316794 534454 317414 569898
rect 316794 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 317414 534454
rect 316794 534134 317414 534218
rect 316794 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 317414 534134
rect 316794 498454 317414 533898
rect 316794 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 317414 498454
rect 316794 498134 317414 498218
rect 316794 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 317414 498134
rect 316794 462454 317414 497898
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 318454 317414 353898
rect 316794 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 317414 318454
rect 316794 318134 317414 318218
rect 316794 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 317414 318134
rect 316794 282454 317414 317898
rect 316794 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 317414 282454
rect 316794 282134 317414 282218
rect 316794 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 317414 282134
rect 316794 246454 317414 281898
rect 316794 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 317414 246454
rect 316794 246134 317414 246218
rect 316794 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 317414 246134
rect 316794 210454 317414 245898
rect 316794 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 317414 210454
rect 316794 210134 317414 210218
rect 316794 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 317414 210134
rect 316794 174454 317414 209898
rect 316794 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 317414 174454
rect 316794 174134 317414 174218
rect 316794 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 317414 174134
rect 316794 138454 317414 173898
rect 316794 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 317414 138454
rect 316794 138134 317414 138218
rect 316794 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 317414 138134
rect 316794 102454 317414 137898
rect 316794 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 317414 102454
rect 316794 102134 317414 102218
rect 316794 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 317414 102134
rect 316794 66454 317414 101898
rect 316794 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 317414 66454
rect 316794 66134 317414 66218
rect 316794 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 317414 66134
rect 316794 30454 317414 65898
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 610954 321914 646398
rect 321294 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 321914 610954
rect 321294 610634 321914 610718
rect 321294 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 321914 610634
rect 321294 574954 321914 610398
rect 321294 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 321914 574954
rect 321294 574634 321914 574718
rect 321294 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 321914 574634
rect 321294 538954 321914 574398
rect 321294 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 321914 538954
rect 321294 538634 321914 538718
rect 321294 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 321914 538634
rect 321294 502954 321914 538398
rect 321294 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 321914 502954
rect 321294 502634 321914 502718
rect 321294 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 321914 502634
rect 321294 466954 321914 502398
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 322954 321914 358398
rect 321294 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 321914 322954
rect 321294 322634 321914 322718
rect 321294 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 321914 322634
rect 321294 286954 321914 322398
rect 321294 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 321914 286954
rect 321294 286634 321914 286718
rect 321294 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 321914 286634
rect 321294 250954 321914 286398
rect 321294 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 321914 250954
rect 321294 250634 321914 250718
rect 321294 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 321914 250634
rect 321294 214954 321914 250398
rect 321294 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 321914 214954
rect 321294 214634 321914 214718
rect 321294 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 321914 214634
rect 321294 178954 321914 214398
rect 321294 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 321914 178954
rect 321294 178634 321914 178718
rect 321294 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 321914 178634
rect 321294 142954 321914 178398
rect 321294 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 321914 142954
rect 321294 142634 321914 142718
rect 321294 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 321914 142634
rect 321294 106954 321914 142398
rect 321294 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 321914 106954
rect 321294 106634 321914 106718
rect 321294 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 321914 106634
rect 321294 70954 321914 106398
rect 321294 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 321914 70954
rect 321294 70634 321914 70718
rect 321294 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 321914 70634
rect 321294 34954 321914 70398
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 331954 330914 367398
rect 330294 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 330914 331954
rect 330294 331634 330914 331718
rect 330294 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 330914 331634
rect 330294 295954 330914 331398
rect 330294 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 330914 295954
rect 330294 295634 330914 295718
rect 330294 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 330914 295634
rect 330294 259954 330914 295398
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 187954 330914 223398
rect 330294 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 330914 187954
rect 330294 187634 330914 187718
rect 330294 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 330914 187634
rect 330294 151954 330914 187398
rect 330294 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 330914 151954
rect 330294 151634 330914 151718
rect 330294 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 330914 151634
rect 330294 115954 330914 151398
rect 330294 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 330914 115954
rect 330294 115634 330914 115718
rect 330294 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 330914 115634
rect 330294 79954 330914 115398
rect 330294 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 330914 79954
rect 330294 79634 330914 79718
rect 330294 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 330914 79634
rect 330294 43954 330914 79398
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 300454 335414 335898
rect 334794 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 335414 300454
rect 334794 300134 335414 300218
rect 334794 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 335414 300134
rect 334794 264454 335414 299898
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 192454 335414 227898
rect 334794 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 335414 192454
rect 334794 192134 335414 192218
rect 334794 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 335414 192134
rect 334794 156454 335414 191898
rect 334794 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 335414 156454
rect 334794 156134 335414 156218
rect 334794 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 335414 156134
rect 334794 120454 335414 155898
rect 334794 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 335414 120454
rect 334794 120134 335414 120218
rect 334794 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 335414 120134
rect 334794 84454 335414 119898
rect 334794 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 335414 84454
rect 334794 84134 335414 84218
rect 334794 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 335414 84134
rect 334794 48454 335414 83898
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 304954 339914 340398
rect 339294 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 339914 304954
rect 339294 304634 339914 304718
rect 339294 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 339914 304634
rect 339294 268954 339914 304398
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 196954 339914 232398
rect 339294 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 339914 196954
rect 339294 196634 339914 196718
rect 339294 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 339914 196634
rect 339294 160954 339914 196398
rect 339294 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 339914 160954
rect 339294 160634 339914 160718
rect 339294 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 339914 160634
rect 339294 124954 339914 160398
rect 339294 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 339914 124954
rect 339294 124634 339914 124718
rect 339294 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 339914 124634
rect 339294 88954 339914 124398
rect 339294 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 339914 88954
rect 339294 88634 339914 88718
rect 339294 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 339914 88634
rect 339294 52954 339914 88398
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 313954 348914 349398
rect 348294 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 348914 313954
rect 348294 313634 348914 313718
rect 348294 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 348914 313634
rect 348294 277954 348914 313398
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 352794 606454 353414 641898
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 318454 353414 353898
rect 352794 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 353414 318454
rect 352794 318134 353414 318218
rect 352794 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 353414 318134
rect 352794 282454 353414 317898
rect 352794 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 353414 282454
rect 352794 282134 353414 282218
rect 352794 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 353414 282134
rect 352794 246454 353414 281898
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 610954 357914 646398
rect 357294 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 357914 610954
rect 357294 610634 357914 610718
rect 357294 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 357914 610634
rect 357294 574954 357914 610398
rect 357294 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 357914 574954
rect 357294 574634 357914 574718
rect 357294 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 357914 574634
rect 357294 538954 357914 574398
rect 357294 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 357914 538954
rect 357294 538634 357914 538718
rect 357294 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 357914 538634
rect 357294 502954 357914 538398
rect 357294 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 357914 502954
rect 357294 502634 357914 502718
rect 357294 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 357914 502634
rect 357294 466954 357914 502398
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 619954 366914 655398
rect 366294 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 366914 619954
rect 366294 619634 366914 619718
rect 366294 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 366914 619634
rect 366294 583954 366914 619398
rect 366294 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 366914 583954
rect 366294 583634 366914 583718
rect 366294 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 366914 583634
rect 366294 547954 366914 583398
rect 366294 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 366914 547954
rect 366294 547634 366914 547718
rect 366294 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 366914 547634
rect 366294 511954 366914 547398
rect 366294 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 366914 511954
rect 366294 511634 366914 511718
rect 366294 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 366914 511634
rect 366294 475954 366914 511398
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 624454 371414 659898
rect 370794 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 371414 624454
rect 370794 624134 371414 624218
rect 370794 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 371414 624134
rect 370794 588454 371414 623898
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552454 371414 587898
rect 370794 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 371414 552454
rect 370794 552134 371414 552218
rect 370794 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 371414 552134
rect 370794 516454 371414 551898
rect 370794 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 371414 516454
rect 370794 516134 371414 516218
rect 370794 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 371414 516134
rect 370794 480454 371414 515898
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 628954 375914 664398
rect 375294 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 375914 628954
rect 375294 628634 375914 628718
rect 375294 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 375914 628634
rect 375294 592954 375914 628398
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 375294 556954 375914 592398
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 520954 375914 556398
rect 375294 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 375914 520954
rect 375294 520634 375914 520718
rect 375294 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 375914 520634
rect 375294 484954 375914 520398
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 637954 384914 673398
rect 384294 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 384914 637954
rect 384294 637634 384914 637718
rect 384294 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 384914 637634
rect 384294 601954 384914 637398
rect 384294 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 384914 601954
rect 384294 601634 384914 601718
rect 384294 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 384914 601634
rect 384294 565954 384914 601398
rect 384294 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 384914 565954
rect 384294 565634 384914 565718
rect 384294 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 384914 565634
rect 384294 529954 384914 565398
rect 384294 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 384914 529954
rect 384294 529634 384914 529718
rect 384294 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 384914 529634
rect 384294 493954 384914 529398
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642454 389414 677898
rect 388794 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 389414 642454
rect 388794 642134 389414 642218
rect 388794 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 389414 642134
rect 388794 606454 389414 641898
rect 388794 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 389414 606454
rect 388794 606134 389414 606218
rect 388794 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 389414 606134
rect 388794 570454 389414 605898
rect 388794 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 389414 570454
rect 388794 570134 389414 570218
rect 388794 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 389414 570134
rect 388794 534454 389414 569898
rect 388794 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 389414 534454
rect 388794 534134 389414 534218
rect 388794 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 389414 534134
rect 388794 498454 389414 533898
rect 388794 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 389414 498454
rect 388794 498134 389414 498218
rect 388794 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 389414 498134
rect 388794 462454 389414 497898
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 610954 393914 646398
rect 393294 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 393914 610954
rect 393294 610634 393914 610718
rect 393294 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 393914 610634
rect 393294 574954 393914 610398
rect 393294 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 393914 574954
rect 393294 574634 393914 574718
rect 393294 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 393914 574634
rect 393294 538954 393914 574398
rect 393294 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 393914 538954
rect 393294 538634 393914 538718
rect 393294 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 393914 538634
rect 393294 502954 393914 538398
rect 393294 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 393914 502954
rect 393294 502634 393914 502718
rect 393294 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 393914 502634
rect 393294 466954 393914 502398
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 402294 655954 402914 691398
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 619954 402914 655398
rect 402294 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 402914 619954
rect 402294 619634 402914 619718
rect 402294 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 402914 619634
rect 402294 583954 402914 619398
rect 402294 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 402914 583954
rect 402294 583634 402914 583718
rect 402294 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 402914 583634
rect 402294 547954 402914 583398
rect 402294 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 402914 547954
rect 402294 547634 402914 547718
rect 402294 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 402914 547634
rect 402294 511954 402914 547398
rect 402294 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 402914 511954
rect 402294 511634 402914 511718
rect 402294 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 402914 511634
rect 402294 475954 402914 511398
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 624454 479414 659898
rect 478794 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 479414 624454
rect 478794 624134 479414 624218
rect 478794 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 479414 624134
rect 478794 588454 479414 623898
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 516454 479414 551898
rect 478794 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 479414 516454
rect 478794 516134 479414 516218
rect 478794 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 479414 516134
rect 478794 480454 479414 515898
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 628954 483914 664398
rect 483294 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 483914 628954
rect 483294 628634 483914 628718
rect 483294 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 483914 628634
rect 483294 592954 483914 628398
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 520954 483914 556398
rect 483294 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 483914 520954
rect 483294 520634 483914 520718
rect 483294 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 483914 520634
rect 483294 484954 483914 520398
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 492294 637954 492914 673398
rect 492294 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 492914 637954
rect 492294 637634 492914 637718
rect 492294 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 492914 637634
rect 492294 601954 492914 637398
rect 492294 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 492914 601954
rect 492294 601634 492914 601718
rect 492294 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 492914 601634
rect 492294 565954 492914 601398
rect 492294 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 492914 565954
rect 492294 565634 492914 565718
rect 492294 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 492914 565634
rect 492294 529954 492914 565398
rect 492294 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 492914 529954
rect 492294 529634 492914 529718
rect 492294 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 492914 529634
rect 492294 493954 492914 529398
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642454 497414 677898
rect 496794 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 497414 642454
rect 496794 642134 497414 642218
rect 496794 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 497414 642134
rect 496794 606454 497414 641898
rect 496794 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 497414 606454
rect 496794 606134 497414 606218
rect 496794 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 497414 606134
rect 496794 570454 497414 605898
rect 496794 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 497414 570454
rect 496794 570134 497414 570218
rect 496794 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 497414 570134
rect 496794 534454 497414 569898
rect 496794 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 497414 534454
rect 496794 534134 497414 534218
rect 496794 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 497414 534134
rect 496794 498454 497414 533898
rect 496794 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 497414 498454
rect 496794 498134 497414 498218
rect 496794 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 497414 498134
rect 496794 462454 497414 497898
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 610954 501914 646398
rect 501294 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 501914 610954
rect 501294 610634 501914 610718
rect 501294 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 501914 610634
rect 501294 574954 501914 610398
rect 501294 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 501914 574954
rect 501294 574634 501914 574718
rect 501294 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 501914 574634
rect 501294 538954 501914 574398
rect 501294 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 501914 538954
rect 501294 538634 501914 538718
rect 501294 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 501914 538634
rect 501294 502954 501914 538398
rect 501294 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 501914 502954
rect 501294 502634 501914 502718
rect 501294 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 501914 502634
rect 501294 466954 501914 502398
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 619954 510914 655398
rect 510294 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 510914 619954
rect 510294 619634 510914 619718
rect 510294 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 510914 619634
rect 510294 583954 510914 619398
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 510294 511954 510914 547398
rect 510294 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 510914 511954
rect 510294 511634 510914 511718
rect 510294 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 510914 511634
rect 510294 475954 510914 511398
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 624454 515414 659898
rect 514794 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 515414 624454
rect 514794 624134 515414 624218
rect 514794 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 515414 624134
rect 514794 588454 515414 623898
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 516454 515414 551898
rect 514794 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 515414 516454
rect 514794 516134 515414 516218
rect 514794 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 515414 516134
rect 514794 480454 515414 515898
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 514794 -2266 515414 11898
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 628954 519914 664398
rect 519294 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 519914 628954
rect 519294 628634 519914 628718
rect 519294 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 519914 628634
rect 519294 592954 519914 628398
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 520954 519914 556398
rect 519294 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 519914 520954
rect 519294 520634 519914 520718
rect 519294 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 519914 520634
rect 519294 484954 519914 520398
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 519294 -3226 519914 16398
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 580211 697236 580277 697237
rect 580211 697172 580212 697236
rect 580276 697172 580277 697236
rect 580211 697171 580277 697172
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 580214 79389 580274 697171
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 580395 644060 580461 644061
rect 580395 643996 580396 644060
rect 580460 643996 580461 644060
rect 580395 643995 580461 643996
rect 580398 82381 580458 643995
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 580395 82380 580461 82381
rect 580395 82316 580396 82380
rect 580460 82316 580461 82380
rect 580395 82315 580461 82316
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 580211 79388 580277 79389
rect 580211 79324 580212 79388
rect 580276 79324 580277 79388
rect 580211 79323 580277 79324
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 51326 628718 51562 628954
rect 51646 628718 51882 628954
rect 51326 628398 51562 628634
rect 51646 628398 51882 628634
rect 51326 592718 51562 592954
rect 51646 592718 51882 592954
rect 51326 592398 51562 592634
rect 51646 592398 51882 592634
rect 51326 556718 51562 556954
rect 51646 556718 51882 556954
rect 51326 556398 51562 556634
rect 51646 556398 51882 556634
rect 51326 520718 51562 520954
rect 51646 520718 51882 520954
rect 51326 520398 51562 520634
rect 51646 520398 51882 520634
rect 51326 484718 51562 484954
rect 51646 484718 51882 484954
rect 51326 484398 51562 484634
rect 51646 484398 51882 484634
rect 51326 448718 51562 448954
rect 51646 448718 51882 448954
rect 51326 448398 51562 448634
rect 51646 448398 51882 448634
rect 51326 412718 51562 412954
rect 51646 412718 51882 412954
rect 51326 412398 51562 412634
rect 51646 412398 51882 412634
rect 51326 376718 51562 376954
rect 51646 376718 51882 376954
rect 51326 376398 51562 376634
rect 51646 376398 51882 376634
rect 51326 340718 51562 340954
rect 51646 340718 51882 340954
rect 51326 340398 51562 340634
rect 51646 340398 51882 340634
rect 51326 304718 51562 304954
rect 51646 304718 51882 304954
rect 51326 304398 51562 304634
rect 51646 304398 51882 304634
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 60326 637718 60562 637954
rect 60646 637718 60882 637954
rect 60326 637398 60562 637634
rect 60646 637398 60882 637634
rect 60326 601718 60562 601954
rect 60646 601718 60882 601954
rect 60326 601398 60562 601634
rect 60646 601398 60882 601634
rect 60326 565718 60562 565954
rect 60646 565718 60882 565954
rect 60326 565398 60562 565634
rect 60646 565398 60882 565634
rect 60326 529718 60562 529954
rect 60646 529718 60882 529954
rect 60326 529398 60562 529634
rect 60646 529398 60882 529634
rect 60326 493718 60562 493954
rect 60646 493718 60882 493954
rect 60326 493398 60562 493634
rect 60646 493398 60882 493634
rect 60326 457718 60562 457954
rect 60646 457718 60882 457954
rect 60326 457398 60562 457634
rect 60646 457398 60882 457634
rect 60326 421718 60562 421954
rect 60646 421718 60882 421954
rect 60326 421398 60562 421634
rect 60646 421398 60882 421634
rect 60326 385718 60562 385954
rect 60646 385718 60882 385954
rect 60326 385398 60562 385634
rect 60646 385398 60882 385634
rect 60326 349718 60562 349954
rect 60646 349718 60882 349954
rect 60326 349398 60562 349634
rect 60646 349398 60882 349634
rect 60326 313718 60562 313954
rect 60646 313718 60882 313954
rect 60326 313398 60562 313634
rect 60646 313398 60882 313634
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 60326 205718 60562 205954
rect 60646 205718 60882 205954
rect 60326 205398 60562 205634
rect 60646 205398 60882 205634
rect 60326 169718 60562 169954
rect 60646 169718 60882 169954
rect 60326 169398 60562 169634
rect 60646 169398 60882 169634
rect 60326 133718 60562 133954
rect 60646 133718 60882 133954
rect 60326 133398 60562 133634
rect 60646 133398 60882 133634
rect 60326 97718 60562 97954
rect 60646 97718 60882 97954
rect 60326 97398 60562 97634
rect 60646 97398 60882 97634
rect 60326 61718 60562 61954
rect 60646 61718 60882 61954
rect 60326 61398 60562 61634
rect 60646 61398 60882 61634
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 64826 642218 65062 642454
rect 65146 642218 65382 642454
rect 64826 641898 65062 642134
rect 65146 641898 65382 642134
rect 64826 606218 65062 606454
rect 65146 606218 65382 606454
rect 64826 605898 65062 606134
rect 65146 605898 65382 606134
rect 64826 570218 65062 570454
rect 65146 570218 65382 570454
rect 64826 569898 65062 570134
rect 65146 569898 65382 570134
rect 64826 534218 65062 534454
rect 65146 534218 65382 534454
rect 64826 533898 65062 534134
rect 65146 533898 65382 534134
rect 64826 498218 65062 498454
rect 65146 498218 65382 498454
rect 64826 497898 65062 498134
rect 65146 497898 65382 498134
rect 64826 462218 65062 462454
rect 65146 462218 65382 462454
rect 64826 461898 65062 462134
rect 65146 461898 65382 462134
rect 64826 426218 65062 426454
rect 65146 426218 65382 426454
rect 64826 425898 65062 426134
rect 65146 425898 65382 426134
rect 64826 390218 65062 390454
rect 65146 390218 65382 390454
rect 64826 389898 65062 390134
rect 65146 389898 65382 390134
rect 64826 354218 65062 354454
rect 65146 354218 65382 354454
rect 64826 353898 65062 354134
rect 65146 353898 65382 354134
rect 64826 318218 65062 318454
rect 65146 318218 65382 318454
rect 64826 317898 65062 318134
rect 65146 317898 65382 318134
rect 64826 282218 65062 282454
rect 65146 282218 65382 282454
rect 64826 281898 65062 282134
rect 65146 281898 65382 282134
rect 64826 246218 65062 246454
rect 65146 246218 65382 246454
rect 64826 245898 65062 246134
rect 65146 245898 65382 246134
rect 64826 210218 65062 210454
rect 65146 210218 65382 210454
rect 64826 209898 65062 210134
rect 65146 209898 65382 210134
rect 64826 174218 65062 174454
rect 65146 174218 65382 174454
rect 64826 173898 65062 174134
rect 65146 173898 65382 174134
rect 64826 138218 65062 138454
rect 65146 138218 65382 138454
rect 64826 137898 65062 138134
rect 65146 137898 65382 138134
rect 64826 102218 65062 102454
rect 65146 102218 65382 102454
rect 64826 101898 65062 102134
rect 65146 101898 65382 102134
rect 64826 66218 65062 66454
rect 65146 66218 65382 66454
rect 64826 65898 65062 66134
rect 65146 65898 65382 66134
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 69326 646718 69562 646954
rect 69646 646718 69882 646954
rect 69326 646398 69562 646634
rect 69646 646398 69882 646634
rect 69326 610718 69562 610954
rect 69646 610718 69882 610954
rect 69326 610398 69562 610634
rect 69646 610398 69882 610634
rect 69326 574718 69562 574954
rect 69646 574718 69882 574954
rect 69326 574398 69562 574634
rect 69646 574398 69882 574634
rect 69326 538718 69562 538954
rect 69646 538718 69882 538954
rect 69326 538398 69562 538634
rect 69646 538398 69882 538634
rect 69326 502718 69562 502954
rect 69646 502718 69882 502954
rect 69326 502398 69562 502634
rect 69646 502398 69882 502634
rect 69326 466718 69562 466954
rect 69646 466718 69882 466954
rect 69326 466398 69562 466634
rect 69646 466398 69882 466634
rect 69326 430718 69562 430954
rect 69646 430718 69882 430954
rect 69326 430398 69562 430634
rect 69646 430398 69882 430634
rect 69326 394718 69562 394954
rect 69646 394718 69882 394954
rect 69326 394398 69562 394634
rect 69646 394398 69882 394634
rect 69326 358718 69562 358954
rect 69646 358718 69882 358954
rect 69326 358398 69562 358634
rect 69646 358398 69882 358634
rect 69326 322718 69562 322954
rect 69646 322718 69882 322954
rect 69326 322398 69562 322634
rect 69646 322398 69882 322634
rect 69326 286718 69562 286954
rect 69646 286718 69882 286954
rect 69326 286398 69562 286634
rect 69646 286398 69882 286634
rect 69326 250718 69562 250954
rect 69646 250718 69882 250954
rect 69326 250398 69562 250634
rect 69646 250398 69882 250634
rect 69326 214718 69562 214954
rect 69646 214718 69882 214954
rect 69326 214398 69562 214634
rect 69646 214398 69882 214634
rect 69326 178718 69562 178954
rect 69646 178718 69882 178954
rect 69326 178398 69562 178634
rect 69646 178398 69882 178634
rect 69326 142718 69562 142954
rect 69646 142718 69882 142954
rect 69326 142398 69562 142634
rect 69646 142398 69882 142634
rect 69326 106718 69562 106954
rect 69646 106718 69882 106954
rect 69326 106398 69562 106634
rect 69646 106398 69882 106634
rect 69326 70718 69562 70954
rect 69646 70718 69882 70954
rect 69326 70398 69562 70634
rect 69646 70398 69882 70634
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 78326 655718 78562 655954
rect 78646 655718 78882 655954
rect 78326 655398 78562 655634
rect 78646 655398 78882 655634
rect 78326 619718 78562 619954
rect 78646 619718 78882 619954
rect 78326 619398 78562 619634
rect 78646 619398 78882 619634
rect 78326 583718 78562 583954
rect 78646 583718 78882 583954
rect 78326 583398 78562 583634
rect 78646 583398 78882 583634
rect 78326 547718 78562 547954
rect 78646 547718 78882 547954
rect 78326 547398 78562 547634
rect 78646 547398 78882 547634
rect 78326 511718 78562 511954
rect 78646 511718 78882 511954
rect 78326 511398 78562 511634
rect 78646 511398 78882 511634
rect 78326 475718 78562 475954
rect 78646 475718 78882 475954
rect 78326 475398 78562 475634
rect 78646 475398 78882 475634
rect 78326 439718 78562 439954
rect 78646 439718 78882 439954
rect 78326 439398 78562 439634
rect 78646 439398 78882 439634
rect 78326 403718 78562 403954
rect 78646 403718 78882 403954
rect 78326 403398 78562 403634
rect 78646 403398 78882 403634
rect 78326 367718 78562 367954
rect 78646 367718 78882 367954
rect 78326 367398 78562 367634
rect 78646 367398 78882 367634
rect 78326 331718 78562 331954
rect 78646 331718 78882 331954
rect 78326 331398 78562 331634
rect 78646 331398 78882 331634
rect 78326 295718 78562 295954
rect 78646 295718 78882 295954
rect 78326 295398 78562 295634
rect 78646 295398 78882 295634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 78326 187718 78562 187954
rect 78646 187718 78882 187954
rect 78326 187398 78562 187634
rect 78646 187398 78882 187634
rect 78326 151718 78562 151954
rect 78646 151718 78882 151954
rect 78326 151398 78562 151634
rect 78646 151398 78882 151634
rect 78326 115718 78562 115954
rect 78646 115718 78882 115954
rect 78326 115398 78562 115634
rect 78646 115398 78882 115634
rect 78326 79718 78562 79954
rect 78646 79718 78882 79954
rect 78326 79398 78562 79634
rect 78646 79398 78882 79634
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 82826 660218 83062 660454
rect 83146 660218 83382 660454
rect 82826 659898 83062 660134
rect 83146 659898 83382 660134
rect 82826 624218 83062 624454
rect 83146 624218 83382 624454
rect 82826 623898 83062 624134
rect 83146 623898 83382 624134
rect 82826 588218 83062 588454
rect 83146 588218 83382 588454
rect 82826 587898 83062 588134
rect 83146 587898 83382 588134
rect 82826 552218 83062 552454
rect 83146 552218 83382 552454
rect 82826 551898 83062 552134
rect 83146 551898 83382 552134
rect 82826 516218 83062 516454
rect 83146 516218 83382 516454
rect 82826 515898 83062 516134
rect 83146 515898 83382 516134
rect 82826 480218 83062 480454
rect 83146 480218 83382 480454
rect 82826 479898 83062 480134
rect 83146 479898 83382 480134
rect 82826 444218 83062 444454
rect 83146 444218 83382 444454
rect 82826 443898 83062 444134
rect 83146 443898 83382 444134
rect 82826 408218 83062 408454
rect 83146 408218 83382 408454
rect 82826 407898 83062 408134
rect 83146 407898 83382 408134
rect 82826 372218 83062 372454
rect 83146 372218 83382 372454
rect 82826 371898 83062 372134
rect 83146 371898 83382 372134
rect 82826 336218 83062 336454
rect 83146 336218 83382 336454
rect 82826 335898 83062 336134
rect 83146 335898 83382 336134
rect 82826 300218 83062 300454
rect 83146 300218 83382 300454
rect 82826 299898 83062 300134
rect 83146 299898 83382 300134
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 82826 192218 83062 192454
rect 83146 192218 83382 192454
rect 82826 191898 83062 192134
rect 83146 191898 83382 192134
rect 82826 156218 83062 156454
rect 83146 156218 83382 156454
rect 82826 155898 83062 156134
rect 83146 155898 83382 156134
rect 82826 120218 83062 120454
rect 83146 120218 83382 120454
rect 82826 119898 83062 120134
rect 83146 119898 83382 120134
rect 82826 84218 83062 84454
rect 83146 84218 83382 84454
rect 82826 83898 83062 84134
rect 83146 83898 83382 84134
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 87326 628718 87562 628954
rect 87646 628718 87882 628954
rect 87326 628398 87562 628634
rect 87646 628398 87882 628634
rect 87326 592718 87562 592954
rect 87646 592718 87882 592954
rect 87326 592398 87562 592634
rect 87646 592398 87882 592634
rect 87326 556718 87562 556954
rect 87646 556718 87882 556954
rect 87326 556398 87562 556634
rect 87646 556398 87882 556634
rect 87326 520718 87562 520954
rect 87646 520718 87882 520954
rect 87326 520398 87562 520634
rect 87646 520398 87882 520634
rect 87326 484718 87562 484954
rect 87646 484718 87882 484954
rect 87326 484398 87562 484634
rect 87646 484398 87882 484634
rect 87326 448718 87562 448954
rect 87646 448718 87882 448954
rect 87326 448398 87562 448634
rect 87646 448398 87882 448634
rect 87326 412718 87562 412954
rect 87646 412718 87882 412954
rect 87326 412398 87562 412634
rect 87646 412398 87882 412634
rect 87326 376718 87562 376954
rect 87646 376718 87882 376954
rect 87326 376398 87562 376634
rect 87646 376398 87882 376634
rect 87326 340718 87562 340954
rect 87646 340718 87882 340954
rect 87326 340398 87562 340634
rect 87646 340398 87882 340634
rect 87326 304718 87562 304954
rect 87646 304718 87882 304954
rect 87326 304398 87562 304634
rect 87646 304398 87882 304634
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 87326 196718 87562 196954
rect 87646 196718 87882 196954
rect 87326 196398 87562 196634
rect 87646 196398 87882 196634
rect 87326 160718 87562 160954
rect 87646 160718 87882 160954
rect 87326 160398 87562 160634
rect 87646 160398 87882 160634
rect 87326 124718 87562 124954
rect 87646 124718 87882 124954
rect 87326 124398 87562 124634
rect 87646 124398 87882 124634
rect 87326 88718 87562 88954
rect 87646 88718 87882 88954
rect 87326 88398 87562 88634
rect 87646 88398 87882 88634
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 96326 637718 96562 637954
rect 96646 637718 96882 637954
rect 96326 637398 96562 637634
rect 96646 637398 96882 637634
rect 96326 601718 96562 601954
rect 96646 601718 96882 601954
rect 96326 601398 96562 601634
rect 96646 601398 96882 601634
rect 96326 565718 96562 565954
rect 96646 565718 96882 565954
rect 96326 565398 96562 565634
rect 96646 565398 96882 565634
rect 96326 529718 96562 529954
rect 96646 529718 96882 529954
rect 96326 529398 96562 529634
rect 96646 529398 96882 529634
rect 96326 493718 96562 493954
rect 96646 493718 96882 493954
rect 96326 493398 96562 493634
rect 96646 493398 96882 493634
rect 96326 457718 96562 457954
rect 96646 457718 96882 457954
rect 96326 457398 96562 457634
rect 96646 457398 96882 457634
rect 96326 421718 96562 421954
rect 96646 421718 96882 421954
rect 96326 421398 96562 421634
rect 96646 421398 96882 421634
rect 96326 385718 96562 385954
rect 96646 385718 96882 385954
rect 96326 385398 96562 385634
rect 96646 385398 96882 385634
rect 96326 349718 96562 349954
rect 96646 349718 96882 349954
rect 96326 349398 96562 349634
rect 96646 349398 96882 349634
rect 96326 313718 96562 313954
rect 96646 313718 96882 313954
rect 96326 313398 96562 313634
rect 96646 313398 96882 313634
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 96326 205718 96562 205954
rect 96646 205718 96882 205954
rect 96326 205398 96562 205634
rect 96646 205398 96882 205634
rect 96326 169718 96562 169954
rect 96646 169718 96882 169954
rect 96326 169398 96562 169634
rect 96646 169398 96882 169634
rect 96326 133718 96562 133954
rect 96646 133718 96882 133954
rect 96326 133398 96562 133634
rect 96646 133398 96882 133634
rect 96326 97718 96562 97954
rect 96646 97718 96882 97954
rect 96326 97398 96562 97634
rect 96646 97398 96882 97634
rect 96326 61718 96562 61954
rect 96646 61718 96882 61954
rect 96326 61398 96562 61634
rect 96646 61398 96882 61634
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 100826 642218 101062 642454
rect 101146 642218 101382 642454
rect 100826 641898 101062 642134
rect 101146 641898 101382 642134
rect 100826 606218 101062 606454
rect 101146 606218 101382 606454
rect 100826 605898 101062 606134
rect 101146 605898 101382 606134
rect 100826 570218 101062 570454
rect 101146 570218 101382 570454
rect 100826 569898 101062 570134
rect 101146 569898 101382 570134
rect 100826 534218 101062 534454
rect 101146 534218 101382 534454
rect 100826 533898 101062 534134
rect 101146 533898 101382 534134
rect 100826 498218 101062 498454
rect 101146 498218 101382 498454
rect 100826 497898 101062 498134
rect 101146 497898 101382 498134
rect 100826 462218 101062 462454
rect 101146 462218 101382 462454
rect 100826 461898 101062 462134
rect 101146 461898 101382 462134
rect 100826 426218 101062 426454
rect 101146 426218 101382 426454
rect 100826 425898 101062 426134
rect 101146 425898 101382 426134
rect 100826 390218 101062 390454
rect 101146 390218 101382 390454
rect 100826 389898 101062 390134
rect 101146 389898 101382 390134
rect 100826 354218 101062 354454
rect 101146 354218 101382 354454
rect 100826 353898 101062 354134
rect 101146 353898 101382 354134
rect 100826 318218 101062 318454
rect 101146 318218 101382 318454
rect 100826 317898 101062 318134
rect 101146 317898 101382 318134
rect 100826 282218 101062 282454
rect 101146 282218 101382 282454
rect 100826 281898 101062 282134
rect 101146 281898 101382 282134
rect 100826 246218 101062 246454
rect 101146 246218 101382 246454
rect 100826 245898 101062 246134
rect 101146 245898 101382 246134
rect 100826 210218 101062 210454
rect 101146 210218 101382 210454
rect 100826 209898 101062 210134
rect 101146 209898 101382 210134
rect 100826 174218 101062 174454
rect 101146 174218 101382 174454
rect 100826 173898 101062 174134
rect 101146 173898 101382 174134
rect 100826 138218 101062 138454
rect 101146 138218 101382 138454
rect 100826 137898 101062 138134
rect 101146 137898 101382 138134
rect 100826 102218 101062 102454
rect 101146 102218 101382 102454
rect 100826 101898 101062 102134
rect 101146 101898 101382 102134
rect 100826 66218 101062 66454
rect 101146 66218 101382 66454
rect 100826 65898 101062 66134
rect 101146 65898 101382 66134
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 105326 646718 105562 646954
rect 105646 646718 105882 646954
rect 105326 646398 105562 646634
rect 105646 646398 105882 646634
rect 105326 610718 105562 610954
rect 105646 610718 105882 610954
rect 105326 610398 105562 610634
rect 105646 610398 105882 610634
rect 105326 574718 105562 574954
rect 105646 574718 105882 574954
rect 105326 574398 105562 574634
rect 105646 574398 105882 574634
rect 105326 538718 105562 538954
rect 105646 538718 105882 538954
rect 105326 538398 105562 538634
rect 105646 538398 105882 538634
rect 105326 502718 105562 502954
rect 105646 502718 105882 502954
rect 105326 502398 105562 502634
rect 105646 502398 105882 502634
rect 105326 466718 105562 466954
rect 105646 466718 105882 466954
rect 105326 466398 105562 466634
rect 105646 466398 105882 466634
rect 105326 430718 105562 430954
rect 105646 430718 105882 430954
rect 105326 430398 105562 430634
rect 105646 430398 105882 430634
rect 105326 394718 105562 394954
rect 105646 394718 105882 394954
rect 105326 394398 105562 394634
rect 105646 394398 105882 394634
rect 105326 358718 105562 358954
rect 105646 358718 105882 358954
rect 105326 358398 105562 358634
rect 105646 358398 105882 358634
rect 105326 322718 105562 322954
rect 105646 322718 105882 322954
rect 105326 322398 105562 322634
rect 105646 322398 105882 322634
rect 105326 286718 105562 286954
rect 105646 286718 105882 286954
rect 105326 286398 105562 286634
rect 105646 286398 105882 286634
rect 105326 250718 105562 250954
rect 105646 250718 105882 250954
rect 105326 250398 105562 250634
rect 105646 250398 105882 250634
rect 105326 214718 105562 214954
rect 105646 214718 105882 214954
rect 105326 214398 105562 214634
rect 105646 214398 105882 214634
rect 105326 178718 105562 178954
rect 105646 178718 105882 178954
rect 105326 178398 105562 178634
rect 105646 178398 105882 178634
rect 105326 142718 105562 142954
rect 105646 142718 105882 142954
rect 105326 142398 105562 142634
rect 105646 142398 105882 142634
rect 105326 106718 105562 106954
rect 105646 106718 105882 106954
rect 105326 106398 105562 106634
rect 105646 106398 105882 106634
rect 105326 70718 105562 70954
rect 105646 70718 105882 70954
rect 105326 70398 105562 70634
rect 105646 70398 105882 70634
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 114326 655718 114562 655954
rect 114646 655718 114882 655954
rect 114326 655398 114562 655634
rect 114646 655398 114882 655634
rect 114326 619718 114562 619954
rect 114646 619718 114882 619954
rect 114326 619398 114562 619634
rect 114646 619398 114882 619634
rect 114326 583718 114562 583954
rect 114646 583718 114882 583954
rect 114326 583398 114562 583634
rect 114646 583398 114882 583634
rect 114326 547718 114562 547954
rect 114646 547718 114882 547954
rect 114326 547398 114562 547634
rect 114646 547398 114882 547634
rect 114326 511718 114562 511954
rect 114646 511718 114882 511954
rect 114326 511398 114562 511634
rect 114646 511398 114882 511634
rect 114326 475718 114562 475954
rect 114646 475718 114882 475954
rect 114326 475398 114562 475634
rect 114646 475398 114882 475634
rect 114326 439718 114562 439954
rect 114646 439718 114882 439954
rect 114326 439398 114562 439634
rect 114646 439398 114882 439634
rect 114326 403718 114562 403954
rect 114646 403718 114882 403954
rect 114326 403398 114562 403634
rect 114646 403398 114882 403634
rect 114326 367718 114562 367954
rect 114646 367718 114882 367954
rect 114326 367398 114562 367634
rect 114646 367398 114882 367634
rect 114326 331718 114562 331954
rect 114646 331718 114882 331954
rect 114326 331398 114562 331634
rect 114646 331398 114882 331634
rect 114326 295718 114562 295954
rect 114646 295718 114882 295954
rect 114326 295398 114562 295634
rect 114646 295398 114882 295634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 114326 187718 114562 187954
rect 114646 187718 114882 187954
rect 114326 187398 114562 187634
rect 114646 187398 114882 187634
rect 114326 151718 114562 151954
rect 114646 151718 114882 151954
rect 114326 151398 114562 151634
rect 114646 151398 114882 151634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 118826 660218 119062 660454
rect 119146 660218 119382 660454
rect 118826 659898 119062 660134
rect 119146 659898 119382 660134
rect 118826 624218 119062 624454
rect 119146 624218 119382 624454
rect 118826 623898 119062 624134
rect 119146 623898 119382 624134
rect 118826 588218 119062 588454
rect 119146 588218 119382 588454
rect 118826 587898 119062 588134
rect 119146 587898 119382 588134
rect 118826 552218 119062 552454
rect 119146 552218 119382 552454
rect 118826 551898 119062 552134
rect 119146 551898 119382 552134
rect 118826 516218 119062 516454
rect 119146 516218 119382 516454
rect 118826 515898 119062 516134
rect 119146 515898 119382 516134
rect 118826 480218 119062 480454
rect 119146 480218 119382 480454
rect 118826 479898 119062 480134
rect 119146 479898 119382 480134
rect 118826 444218 119062 444454
rect 119146 444218 119382 444454
rect 118826 443898 119062 444134
rect 119146 443898 119382 444134
rect 118826 408218 119062 408454
rect 119146 408218 119382 408454
rect 118826 407898 119062 408134
rect 119146 407898 119382 408134
rect 118826 372218 119062 372454
rect 119146 372218 119382 372454
rect 118826 371898 119062 372134
rect 119146 371898 119382 372134
rect 118826 336218 119062 336454
rect 119146 336218 119382 336454
rect 118826 335898 119062 336134
rect 119146 335898 119382 336134
rect 118826 300218 119062 300454
rect 119146 300218 119382 300454
rect 118826 299898 119062 300134
rect 119146 299898 119382 300134
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 118826 192218 119062 192454
rect 119146 192218 119382 192454
rect 118826 191898 119062 192134
rect 119146 191898 119382 192134
rect 118826 156218 119062 156454
rect 119146 156218 119382 156454
rect 118826 155898 119062 156134
rect 119146 155898 119382 156134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 123326 628718 123562 628954
rect 123646 628718 123882 628954
rect 123326 628398 123562 628634
rect 123646 628398 123882 628634
rect 123326 592718 123562 592954
rect 123646 592718 123882 592954
rect 123326 592398 123562 592634
rect 123646 592398 123882 592634
rect 123326 556718 123562 556954
rect 123646 556718 123882 556954
rect 123326 556398 123562 556634
rect 123646 556398 123882 556634
rect 123326 520718 123562 520954
rect 123646 520718 123882 520954
rect 123326 520398 123562 520634
rect 123646 520398 123882 520634
rect 123326 484718 123562 484954
rect 123646 484718 123882 484954
rect 123326 484398 123562 484634
rect 123646 484398 123882 484634
rect 123326 448718 123562 448954
rect 123646 448718 123882 448954
rect 123326 448398 123562 448634
rect 123646 448398 123882 448634
rect 123326 412718 123562 412954
rect 123646 412718 123882 412954
rect 123326 412398 123562 412634
rect 123646 412398 123882 412634
rect 123326 376718 123562 376954
rect 123646 376718 123882 376954
rect 123326 376398 123562 376634
rect 123646 376398 123882 376634
rect 123326 340718 123562 340954
rect 123646 340718 123882 340954
rect 123326 340398 123562 340634
rect 123646 340398 123882 340634
rect 123326 304718 123562 304954
rect 123646 304718 123882 304954
rect 123326 304398 123562 304634
rect 123646 304398 123882 304634
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 123326 196718 123562 196954
rect 123646 196718 123882 196954
rect 123326 196398 123562 196634
rect 123646 196398 123882 196634
rect 123326 160718 123562 160954
rect 123646 160718 123882 160954
rect 123326 160398 123562 160634
rect 123646 160398 123882 160634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 132326 637718 132562 637954
rect 132646 637718 132882 637954
rect 132326 637398 132562 637634
rect 132646 637398 132882 637634
rect 132326 601718 132562 601954
rect 132646 601718 132882 601954
rect 132326 601398 132562 601634
rect 132646 601398 132882 601634
rect 132326 565718 132562 565954
rect 132646 565718 132882 565954
rect 132326 565398 132562 565634
rect 132646 565398 132882 565634
rect 132326 529718 132562 529954
rect 132646 529718 132882 529954
rect 132326 529398 132562 529634
rect 132646 529398 132882 529634
rect 132326 493718 132562 493954
rect 132646 493718 132882 493954
rect 132326 493398 132562 493634
rect 132646 493398 132882 493634
rect 132326 457718 132562 457954
rect 132646 457718 132882 457954
rect 132326 457398 132562 457634
rect 132646 457398 132882 457634
rect 132326 421718 132562 421954
rect 132646 421718 132882 421954
rect 132326 421398 132562 421634
rect 132646 421398 132882 421634
rect 132326 385718 132562 385954
rect 132646 385718 132882 385954
rect 132326 385398 132562 385634
rect 132646 385398 132882 385634
rect 132326 349718 132562 349954
rect 132646 349718 132882 349954
rect 132326 349398 132562 349634
rect 132646 349398 132882 349634
rect 132326 313718 132562 313954
rect 132646 313718 132882 313954
rect 132326 313398 132562 313634
rect 132646 313398 132882 313634
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 132326 205718 132562 205954
rect 132646 205718 132882 205954
rect 132326 205398 132562 205634
rect 132646 205398 132882 205634
rect 132326 169718 132562 169954
rect 132646 169718 132882 169954
rect 132326 169398 132562 169634
rect 132646 169398 132882 169634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 136826 642218 137062 642454
rect 137146 642218 137382 642454
rect 136826 641898 137062 642134
rect 137146 641898 137382 642134
rect 136826 606218 137062 606454
rect 137146 606218 137382 606454
rect 136826 605898 137062 606134
rect 137146 605898 137382 606134
rect 136826 570218 137062 570454
rect 137146 570218 137382 570454
rect 136826 569898 137062 570134
rect 137146 569898 137382 570134
rect 136826 534218 137062 534454
rect 137146 534218 137382 534454
rect 136826 533898 137062 534134
rect 137146 533898 137382 534134
rect 136826 498218 137062 498454
rect 137146 498218 137382 498454
rect 136826 497898 137062 498134
rect 137146 497898 137382 498134
rect 136826 462218 137062 462454
rect 137146 462218 137382 462454
rect 136826 461898 137062 462134
rect 137146 461898 137382 462134
rect 136826 426218 137062 426454
rect 137146 426218 137382 426454
rect 136826 425898 137062 426134
rect 137146 425898 137382 426134
rect 136826 390218 137062 390454
rect 137146 390218 137382 390454
rect 136826 389898 137062 390134
rect 137146 389898 137382 390134
rect 136826 354218 137062 354454
rect 137146 354218 137382 354454
rect 136826 353898 137062 354134
rect 137146 353898 137382 354134
rect 136826 318218 137062 318454
rect 137146 318218 137382 318454
rect 136826 317898 137062 318134
rect 137146 317898 137382 318134
rect 136826 282218 137062 282454
rect 137146 282218 137382 282454
rect 136826 281898 137062 282134
rect 137146 281898 137382 282134
rect 136826 246218 137062 246454
rect 137146 246218 137382 246454
rect 136826 245898 137062 246134
rect 137146 245898 137382 246134
rect 136826 210218 137062 210454
rect 137146 210218 137382 210454
rect 136826 209898 137062 210134
rect 137146 209898 137382 210134
rect 136826 174218 137062 174454
rect 137146 174218 137382 174454
rect 136826 173898 137062 174134
rect 137146 173898 137382 174134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 141326 646718 141562 646954
rect 141646 646718 141882 646954
rect 141326 646398 141562 646634
rect 141646 646398 141882 646634
rect 141326 610718 141562 610954
rect 141646 610718 141882 610954
rect 141326 610398 141562 610634
rect 141646 610398 141882 610634
rect 141326 574718 141562 574954
rect 141646 574718 141882 574954
rect 141326 574398 141562 574634
rect 141646 574398 141882 574634
rect 141326 538718 141562 538954
rect 141646 538718 141882 538954
rect 141326 538398 141562 538634
rect 141646 538398 141882 538634
rect 141326 502718 141562 502954
rect 141646 502718 141882 502954
rect 141326 502398 141562 502634
rect 141646 502398 141882 502634
rect 141326 466718 141562 466954
rect 141646 466718 141882 466954
rect 141326 466398 141562 466634
rect 141646 466398 141882 466634
rect 141326 430718 141562 430954
rect 141646 430718 141882 430954
rect 141326 430398 141562 430634
rect 141646 430398 141882 430634
rect 141326 394718 141562 394954
rect 141646 394718 141882 394954
rect 141326 394398 141562 394634
rect 141646 394398 141882 394634
rect 141326 358718 141562 358954
rect 141646 358718 141882 358954
rect 141326 358398 141562 358634
rect 141646 358398 141882 358634
rect 141326 322718 141562 322954
rect 141646 322718 141882 322954
rect 141326 322398 141562 322634
rect 141646 322398 141882 322634
rect 141326 286718 141562 286954
rect 141646 286718 141882 286954
rect 141326 286398 141562 286634
rect 141646 286398 141882 286634
rect 141326 250718 141562 250954
rect 141646 250718 141882 250954
rect 141326 250398 141562 250634
rect 141646 250398 141882 250634
rect 141326 214718 141562 214954
rect 141646 214718 141882 214954
rect 141326 214398 141562 214634
rect 141646 214398 141882 214634
rect 141326 178718 141562 178954
rect 141646 178718 141882 178954
rect 141326 178398 141562 178634
rect 141646 178398 141882 178634
rect 141326 142718 141562 142954
rect 141646 142718 141882 142954
rect 141326 142398 141562 142634
rect 141646 142398 141882 142634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 150326 655718 150562 655954
rect 150646 655718 150882 655954
rect 150326 655398 150562 655634
rect 150646 655398 150882 655634
rect 150326 619718 150562 619954
rect 150646 619718 150882 619954
rect 150326 619398 150562 619634
rect 150646 619398 150882 619634
rect 150326 583718 150562 583954
rect 150646 583718 150882 583954
rect 150326 583398 150562 583634
rect 150646 583398 150882 583634
rect 150326 547718 150562 547954
rect 150646 547718 150882 547954
rect 150326 547398 150562 547634
rect 150646 547398 150882 547634
rect 150326 511718 150562 511954
rect 150646 511718 150882 511954
rect 150326 511398 150562 511634
rect 150646 511398 150882 511634
rect 150326 475718 150562 475954
rect 150646 475718 150882 475954
rect 150326 475398 150562 475634
rect 150646 475398 150882 475634
rect 150326 439718 150562 439954
rect 150646 439718 150882 439954
rect 150326 439398 150562 439634
rect 150646 439398 150882 439634
rect 150326 403718 150562 403954
rect 150646 403718 150882 403954
rect 150326 403398 150562 403634
rect 150646 403398 150882 403634
rect 150326 367718 150562 367954
rect 150646 367718 150882 367954
rect 150326 367398 150562 367634
rect 150646 367398 150882 367634
rect 150326 331718 150562 331954
rect 150646 331718 150882 331954
rect 150326 331398 150562 331634
rect 150646 331398 150882 331634
rect 150326 295718 150562 295954
rect 150646 295718 150882 295954
rect 150326 295398 150562 295634
rect 150646 295398 150882 295634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 150326 187718 150562 187954
rect 150646 187718 150882 187954
rect 150326 187398 150562 187634
rect 150646 187398 150882 187634
rect 150326 151718 150562 151954
rect 150646 151718 150882 151954
rect 150326 151398 150562 151634
rect 150646 151398 150882 151634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 154826 660218 155062 660454
rect 155146 660218 155382 660454
rect 154826 659898 155062 660134
rect 155146 659898 155382 660134
rect 154826 624218 155062 624454
rect 155146 624218 155382 624454
rect 154826 623898 155062 624134
rect 155146 623898 155382 624134
rect 154826 588218 155062 588454
rect 155146 588218 155382 588454
rect 154826 587898 155062 588134
rect 155146 587898 155382 588134
rect 154826 552218 155062 552454
rect 155146 552218 155382 552454
rect 154826 551898 155062 552134
rect 155146 551898 155382 552134
rect 154826 516218 155062 516454
rect 155146 516218 155382 516454
rect 154826 515898 155062 516134
rect 155146 515898 155382 516134
rect 154826 480218 155062 480454
rect 155146 480218 155382 480454
rect 154826 479898 155062 480134
rect 155146 479898 155382 480134
rect 154826 444218 155062 444454
rect 155146 444218 155382 444454
rect 154826 443898 155062 444134
rect 155146 443898 155382 444134
rect 154826 408218 155062 408454
rect 155146 408218 155382 408454
rect 154826 407898 155062 408134
rect 155146 407898 155382 408134
rect 154826 372218 155062 372454
rect 155146 372218 155382 372454
rect 154826 371898 155062 372134
rect 155146 371898 155382 372134
rect 154826 336218 155062 336454
rect 155146 336218 155382 336454
rect 154826 335898 155062 336134
rect 155146 335898 155382 336134
rect 154826 300218 155062 300454
rect 155146 300218 155382 300454
rect 154826 299898 155062 300134
rect 155146 299898 155382 300134
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 154826 192218 155062 192454
rect 155146 192218 155382 192454
rect 154826 191898 155062 192134
rect 155146 191898 155382 192134
rect 154826 156218 155062 156454
rect 155146 156218 155382 156454
rect 154826 155898 155062 156134
rect 155146 155898 155382 156134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 159326 628718 159562 628954
rect 159646 628718 159882 628954
rect 159326 628398 159562 628634
rect 159646 628398 159882 628634
rect 159326 592718 159562 592954
rect 159646 592718 159882 592954
rect 159326 592398 159562 592634
rect 159646 592398 159882 592634
rect 159326 556718 159562 556954
rect 159646 556718 159882 556954
rect 159326 556398 159562 556634
rect 159646 556398 159882 556634
rect 159326 520718 159562 520954
rect 159646 520718 159882 520954
rect 159326 520398 159562 520634
rect 159646 520398 159882 520634
rect 159326 484718 159562 484954
rect 159646 484718 159882 484954
rect 159326 484398 159562 484634
rect 159646 484398 159882 484634
rect 159326 448718 159562 448954
rect 159646 448718 159882 448954
rect 159326 448398 159562 448634
rect 159646 448398 159882 448634
rect 159326 412718 159562 412954
rect 159646 412718 159882 412954
rect 159326 412398 159562 412634
rect 159646 412398 159882 412634
rect 159326 376718 159562 376954
rect 159646 376718 159882 376954
rect 159326 376398 159562 376634
rect 159646 376398 159882 376634
rect 159326 340718 159562 340954
rect 159646 340718 159882 340954
rect 159326 340398 159562 340634
rect 159646 340398 159882 340634
rect 159326 304718 159562 304954
rect 159646 304718 159882 304954
rect 159326 304398 159562 304634
rect 159646 304398 159882 304634
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 159326 196718 159562 196954
rect 159646 196718 159882 196954
rect 159326 196398 159562 196634
rect 159646 196398 159882 196634
rect 159326 160718 159562 160954
rect 159646 160718 159882 160954
rect 159326 160398 159562 160634
rect 159646 160398 159882 160634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 168326 637718 168562 637954
rect 168646 637718 168882 637954
rect 168326 637398 168562 637634
rect 168646 637398 168882 637634
rect 168326 601718 168562 601954
rect 168646 601718 168882 601954
rect 168326 601398 168562 601634
rect 168646 601398 168882 601634
rect 168326 565718 168562 565954
rect 168646 565718 168882 565954
rect 168326 565398 168562 565634
rect 168646 565398 168882 565634
rect 168326 529718 168562 529954
rect 168646 529718 168882 529954
rect 168326 529398 168562 529634
rect 168646 529398 168882 529634
rect 168326 493718 168562 493954
rect 168646 493718 168882 493954
rect 168326 493398 168562 493634
rect 168646 493398 168882 493634
rect 168326 457718 168562 457954
rect 168646 457718 168882 457954
rect 168326 457398 168562 457634
rect 168646 457398 168882 457634
rect 168326 421718 168562 421954
rect 168646 421718 168882 421954
rect 168326 421398 168562 421634
rect 168646 421398 168882 421634
rect 168326 385718 168562 385954
rect 168646 385718 168882 385954
rect 168326 385398 168562 385634
rect 168646 385398 168882 385634
rect 168326 349718 168562 349954
rect 168646 349718 168882 349954
rect 168326 349398 168562 349634
rect 168646 349398 168882 349634
rect 168326 313718 168562 313954
rect 168646 313718 168882 313954
rect 168326 313398 168562 313634
rect 168646 313398 168882 313634
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 168326 205718 168562 205954
rect 168646 205718 168882 205954
rect 168326 205398 168562 205634
rect 168646 205398 168882 205634
rect 168326 169718 168562 169954
rect 168646 169718 168882 169954
rect 168326 169398 168562 169634
rect 168646 169398 168882 169634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 172826 642218 173062 642454
rect 173146 642218 173382 642454
rect 172826 641898 173062 642134
rect 173146 641898 173382 642134
rect 172826 606218 173062 606454
rect 173146 606218 173382 606454
rect 172826 605898 173062 606134
rect 173146 605898 173382 606134
rect 172826 570218 173062 570454
rect 173146 570218 173382 570454
rect 172826 569898 173062 570134
rect 173146 569898 173382 570134
rect 172826 534218 173062 534454
rect 173146 534218 173382 534454
rect 172826 533898 173062 534134
rect 173146 533898 173382 534134
rect 172826 498218 173062 498454
rect 173146 498218 173382 498454
rect 172826 497898 173062 498134
rect 173146 497898 173382 498134
rect 172826 462218 173062 462454
rect 173146 462218 173382 462454
rect 172826 461898 173062 462134
rect 173146 461898 173382 462134
rect 172826 426218 173062 426454
rect 173146 426218 173382 426454
rect 172826 425898 173062 426134
rect 173146 425898 173382 426134
rect 172826 390218 173062 390454
rect 173146 390218 173382 390454
rect 172826 389898 173062 390134
rect 173146 389898 173382 390134
rect 172826 354218 173062 354454
rect 173146 354218 173382 354454
rect 172826 353898 173062 354134
rect 173146 353898 173382 354134
rect 172826 318218 173062 318454
rect 173146 318218 173382 318454
rect 172826 317898 173062 318134
rect 173146 317898 173382 318134
rect 172826 282218 173062 282454
rect 173146 282218 173382 282454
rect 172826 281898 173062 282134
rect 173146 281898 173382 282134
rect 172826 246218 173062 246454
rect 173146 246218 173382 246454
rect 172826 245898 173062 246134
rect 173146 245898 173382 246134
rect 172826 210218 173062 210454
rect 173146 210218 173382 210454
rect 172826 209898 173062 210134
rect 173146 209898 173382 210134
rect 172826 174218 173062 174454
rect 173146 174218 173382 174454
rect 172826 173898 173062 174134
rect 173146 173898 173382 174134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 177326 646718 177562 646954
rect 177646 646718 177882 646954
rect 177326 646398 177562 646634
rect 177646 646398 177882 646634
rect 177326 610718 177562 610954
rect 177646 610718 177882 610954
rect 177326 610398 177562 610634
rect 177646 610398 177882 610634
rect 177326 574718 177562 574954
rect 177646 574718 177882 574954
rect 177326 574398 177562 574634
rect 177646 574398 177882 574634
rect 177326 538718 177562 538954
rect 177646 538718 177882 538954
rect 177326 538398 177562 538634
rect 177646 538398 177882 538634
rect 177326 502718 177562 502954
rect 177646 502718 177882 502954
rect 177326 502398 177562 502634
rect 177646 502398 177882 502634
rect 177326 466718 177562 466954
rect 177646 466718 177882 466954
rect 177326 466398 177562 466634
rect 177646 466398 177882 466634
rect 177326 430718 177562 430954
rect 177646 430718 177882 430954
rect 177326 430398 177562 430634
rect 177646 430398 177882 430634
rect 177326 394718 177562 394954
rect 177646 394718 177882 394954
rect 177326 394398 177562 394634
rect 177646 394398 177882 394634
rect 177326 358718 177562 358954
rect 177646 358718 177882 358954
rect 177326 358398 177562 358634
rect 177646 358398 177882 358634
rect 177326 322718 177562 322954
rect 177646 322718 177882 322954
rect 177326 322398 177562 322634
rect 177646 322398 177882 322634
rect 177326 286718 177562 286954
rect 177646 286718 177882 286954
rect 177326 286398 177562 286634
rect 177646 286398 177882 286634
rect 177326 250718 177562 250954
rect 177646 250718 177882 250954
rect 177326 250398 177562 250634
rect 177646 250398 177882 250634
rect 177326 214718 177562 214954
rect 177646 214718 177882 214954
rect 177326 214398 177562 214634
rect 177646 214398 177882 214634
rect 177326 178718 177562 178954
rect 177646 178718 177882 178954
rect 177326 178398 177562 178634
rect 177646 178398 177882 178634
rect 177326 142718 177562 142954
rect 177646 142718 177882 142954
rect 177326 142398 177562 142634
rect 177646 142398 177882 142634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 186326 655718 186562 655954
rect 186646 655718 186882 655954
rect 186326 655398 186562 655634
rect 186646 655398 186882 655634
rect 186326 619718 186562 619954
rect 186646 619718 186882 619954
rect 186326 619398 186562 619634
rect 186646 619398 186882 619634
rect 186326 583718 186562 583954
rect 186646 583718 186882 583954
rect 186326 583398 186562 583634
rect 186646 583398 186882 583634
rect 186326 547718 186562 547954
rect 186646 547718 186882 547954
rect 186326 547398 186562 547634
rect 186646 547398 186882 547634
rect 186326 511718 186562 511954
rect 186646 511718 186882 511954
rect 186326 511398 186562 511634
rect 186646 511398 186882 511634
rect 186326 475718 186562 475954
rect 186646 475718 186882 475954
rect 186326 475398 186562 475634
rect 186646 475398 186882 475634
rect 186326 439718 186562 439954
rect 186646 439718 186882 439954
rect 186326 439398 186562 439634
rect 186646 439398 186882 439634
rect 186326 403718 186562 403954
rect 186646 403718 186882 403954
rect 186326 403398 186562 403634
rect 186646 403398 186882 403634
rect 186326 367718 186562 367954
rect 186646 367718 186882 367954
rect 186326 367398 186562 367634
rect 186646 367398 186882 367634
rect 186326 331718 186562 331954
rect 186646 331718 186882 331954
rect 186326 331398 186562 331634
rect 186646 331398 186882 331634
rect 186326 295718 186562 295954
rect 186646 295718 186882 295954
rect 186326 295398 186562 295634
rect 186646 295398 186882 295634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 186326 187718 186562 187954
rect 186646 187718 186882 187954
rect 186326 187398 186562 187634
rect 186646 187398 186882 187634
rect 186326 151718 186562 151954
rect 186646 151718 186882 151954
rect 186326 151398 186562 151634
rect 186646 151398 186882 151634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 190826 660218 191062 660454
rect 191146 660218 191382 660454
rect 190826 659898 191062 660134
rect 191146 659898 191382 660134
rect 190826 624218 191062 624454
rect 191146 624218 191382 624454
rect 190826 623898 191062 624134
rect 191146 623898 191382 624134
rect 190826 588218 191062 588454
rect 191146 588218 191382 588454
rect 190826 587898 191062 588134
rect 191146 587898 191382 588134
rect 190826 552218 191062 552454
rect 191146 552218 191382 552454
rect 190826 551898 191062 552134
rect 191146 551898 191382 552134
rect 190826 516218 191062 516454
rect 191146 516218 191382 516454
rect 190826 515898 191062 516134
rect 191146 515898 191382 516134
rect 190826 480218 191062 480454
rect 191146 480218 191382 480454
rect 190826 479898 191062 480134
rect 191146 479898 191382 480134
rect 190826 444218 191062 444454
rect 191146 444218 191382 444454
rect 190826 443898 191062 444134
rect 191146 443898 191382 444134
rect 190826 408218 191062 408454
rect 191146 408218 191382 408454
rect 190826 407898 191062 408134
rect 191146 407898 191382 408134
rect 190826 372218 191062 372454
rect 191146 372218 191382 372454
rect 190826 371898 191062 372134
rect 191146 371898 191382 372134
rect 190826 336218 191062 336454
rect 191146 336218 191382 336454
rect 190826 335898 191062 336134
rect 191146 335898 191382 336134
rect 190826 300218 191062 300454
rect 191146 300218 191382 300454
rect 190826 299898 191062 300134
rect 191146 299898 191382 300134
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 190826 192218 191062 192454
rect 191146 192218 191382 192454
rect 190826 191898 191062 192134
rect 191146 191898 191382 192134
rect 190826 156218 191062 156454
rect 191146 156218 191382 156454
rect 190826 155898 191062 156134
rect 191146 155898 191382 156134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 195326 628718 195562 628954
rect 195646 628718 195882 628954
rect 195326 628398 195562 628634
rect 195646 628398 195882 628634
rect 195326 592718 195562 592954
rect 195646 592718 195882 592954
rect 195326 592398 195562 592634
rect 195646 592398 195882 592634
rect 195326 556718 195562 556954
rect 195646 556718 195882 556954
rect 195326 556398 195562 556634
rect 195646 556398 195882 556634
rect 195326 520718 195562 520954
rect 195646 520718 195882 520954
rect 195326 520398 195562 520634
rect 195646 520398 195882 520634
rect 195326 484718 195562 484954
rect 195646 484718 195882 484954
rect 195326 484398 195562 484634
rect 195646 484398 195882 484634
rect 195326 448718 195562 448954
rect 195646 448718 195882 448954
rect 195326 448398 195562 448634
rect 195646 448398 195882 448634
rect 195326 412718 195562 412954
rect 195646 412718 195882 412954
rect 195326 412398 195562 412634
rect 195646 412398 195882 412634
rect 195326 376718 195562 376954
rect 195646 376718 195882 376954
rect 195326 376398 195562 376634
rect 195646 376398 195882 376634
rect 195326 340718 195562 340954
rect 195646 340718 195882 340954
rect 195326 340398 195562 340634
rect 195646 340398 195882 340634
rect 195326 304718 195562 304954
rect 195646 304718 195882 304954
rect 195326 304398 195562 304634
rect 195646 304398 195882 304634
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 195326 196718 195562 196954
rect 195646 196718 195882 196954
rect 195326 196398 195562 196634
rect 195646 196398 195882 196634
rect 195326 160718 195562 160954
rect 195646 160718 195882 160954
rect 195326 160398 195562 160634
rect 195646 160398 195882 160634
rect 195326 124718 195562 124954
rect 195646 124718 195882 124954
rect 195326 124398 195562 124634
rect 195646 124398 195882 124634
rect 114326 115718 114562 115954
rect 114646 115718 114882 115954
rect 114326 115398 114562 115634
rect 114646 115398 114882 115634
rect 139610 115718 139846 115954
rect 139610 115398 139846 115634
rect 170330 115718 170566 115954
rect 170330 115398 170566 115634
rect 124250 111218 124486 111454
rect 124250 110898 124486 111134
rect 154970 111218 155206 111454
rect 154970 110898 155206 111134
rect 185690 111218 185926 111454
rect 185690 110898 185926 111134
rect 195326 88718 195562 88954
rect 195646 88718 195882 88954
rect 195326 88398 195562 88634
rect 195646 88398 195882 88634
rect 114326 79718 114562 79954
rect 114646 79718 114882 79954
rect 114326 79398 114562 79634
rect 114646 79398 114882 79634
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 132326 61718 132562 61954
rect 132646 61718 132882 61954
rect 132326 61398 132562 61634
rect 132646 61398 132882 61634
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 136826 66218 137062 66454
rect 137146 66218 137382 66454
rect 136826 65898 137062 66134
rect 137146 65898 137382 66134
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 141326 70718 141562 70954
rect 141646 70718 141882 70954
rect 141326 70398 141562 70634
rect 141646 70398 141882 70634
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 168326 61718 168562 61954
rect 168646 61718 168882 61954
rect 168326 61398 168562 61634
rect 168646 61398 168882 61634
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 172826 66218 173062 66454
rect 173146 66218 173382 66454
rect 172826 65898 173062 66134
rect 173146 65898 173382 66134
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 177326 70718 177562 70954
rect 177646 70718 177882 70954
rect 177326 70398 177562 70634
rect 177646 70398 177882 70634
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 204326 637718 204562 637954
rect 204646 637718 204882 637954
rect 204326 637398 204562 637634
rect 204646 637398 204882 637634
rect 204326 601718 204562 601954
rect 204646 601718 204882 601954
rect 204326 601398 204562 601634
rect 204646 601398 204882 601634
rect 204326 565718 204562 565954
rect 204646 565718 204882 565954
rect 204326 565398 204562 565634
rect 204646 565398 204882 565634
rect 204326 529718 204562 529954
rect 204646 529718 204882 529954
rect 204326 529398 204562 529634
rect 204646 529398 204882 529634
rect 204326 493718 204562 493954
rect 204646 493718 204882 493954
rect 204326 493398 204562 493634
rect 204646 493398 204882 493634
rect 204326 457718 204562 457954
rect 204646 457718 204882 457954
rect 204326 457398 204562 457634
rect 204646 457398 204882 457634
rect 204326 421718 204562 421954
rect 204646 421718 204882 421954
rect 204326 421398 204562 421634
rect 204646 421398 204882 421634
rect 204326 385718 204562 385954
rect 204646 385718 204882 385954
rect 204326 385398 204562 385634
rect 204646 385398 204882 385634
rect 204326 349718 204562 349954
rect 204646 349718 204882 349954
rect 204326 349398 204562 349634
rect 204646 349398 204882 349634
rect 204326 313718 204562 313954
rect 204646 313718 204882 313954
rect 204326 313398 204562 313634
rect 204646 313398 204882 313634
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 204326 205718 204562 205954
rect 204646 205718 204882 205954
rect 204326 205398 204562 205634
rect 204646 205398 204882 205634
rect 204326 169718 204562 169954
rect 204646 169718 204882 169954
rect 204326 169398 204562 169634
rect 204646 169398 204882 169634
rect 204326 133718 204562 133954
rect 204646 133718 204882 133954
rect 204326 133398 204562 133634
rect 204646 133398 204882 133634
rect 204326 97718 204562 97954
rect 204646 97718 204882 97954
rect 204326 97398 204562 97634
rect 204646 97398 204882 97634
rect 204326 61718 204562 61954
rect 204646 61718 204882 61954
rect 204326 61398 204562 61634
rect 204646 61398 204882 61634
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 208826 642218 209062 642454
rect 209146 642218 209382 642454
rect 208826 641898 209062 642134
rect 209146 641898 209382 642134
rect 208826 606218 209062 606454
rect 209146 606218 209382 606454
rect 208826 605898 209062 606134
rect 209146 605898 209382 606134
rect 208826 570218 209062 570454
rect 209146 570218 209382 570454
rect 208826 569898 209062 570134
rect 209146 569898 209382 570134
rect 208826 534218 209062 534454
rect 209146 534218 209382 534454
rect 208826 533898 209062 534134
rect 209146 533898 209382 534134
rect 208826 498218 209062 498454
rect 209146 498218 209382 498454
rect 208826 497898 209062 498134
rect 209146 497898 209382 498134
rect 208826 462218 209062 462454
rect 209146 462218 209382 462454
rect 208826 461898 209062 462134
rect 209146 461898 209382 462134
rect 208826 426218 209062 426454
rect 209146 426218 209382 426454
rect 208826 425898 209062 426134
rect 209146 425898 209382 426134
rect 208826 390218 209062 390454
rect 209146 390218 209382 390454
rect 208826 389898 209062 390134
rect 209146 389898 209382 390134
rect 208826 354218 209062 354454
rect 209146 354218 209382 354454
rect 208826 353898 209062 354134
rect 209146 353898 209382 354134
rect 208826 318218 209062 318454
rect 209146 318218 209382 318454
rect 208826 317898 209062 318134
rect 209146 317898 209382 318134
rect 208826 282218 209062 282454
rect 209146 282218 209382 282454
rect 208826 281898 209062 282134
rect 209146 281898 209382 282134
rect 208826 246218 209062 246454
rect 209146 246218 209382 246454
rect 208826 245898 209062 246134
rect 209146 245898 209382 246134
rect 208826 210218 209062 210454
rect 209146 210218 209382 210454
rect 208826 209898 209062 210134
rect 209146 209898 209382 210134
rect 208826 174218 209062 174454
rect 209146 174218 209382 174454
rect 208826 173898 209062 174134
rect 209146 173898 209382 174134
rect 208826 138218 209062 138454
rect 209146 138218 209382 138454
rect 208826 137898 209062 138134
rect 209146 137898 209382 138134
rect 208826 102218 209062 102454
rect 209146 102218 209382 102454
rect 208826 101898 209062 102134
rect 209146 101898 209382 102134
rect 208826 66218 209062 66454
rect 209146 66218 209382 66454
rect 208826 65898 209062 66134
rect 209146 65898 209382 66134
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 213326 646718 213562 646954
rect 213646 646718 213882 646954
rect 213326 646398 213562 646634
rect 213646 646398 213882 646634
rect 213326 610718 213562 610954
rect 213646 610718 213882 610954
rect 213326 610398 213562 610634
rect 213646 610398 213882 610634
rect 213326 574718 213562 574954
rect 213646 574718 213882 574954
rect 213326 574398 213562 574634
rect 213646 574398 213882 574634
rect 213326 538718 213562 538954
rect 213646 538718 213882 538954
rect 213326 538398 213562 538634
rect 213646 538398 213882 538634
rect 213326 502718 213562 502954
rect 213646 502718 213882 502954
rect 213326 502398 213562 502634
rect 213646 502398 213882 502634
rect 213326 466718 213562 466954
rect 213646 466718 213882 466954
rect 213326 466398 213562 466634
rect 213646 466398 213882 466634
rect 213326 430718 213562 430954
rect 213646 430718 213882 430954
rect 213326 430398 213562 430634
rect 213646 430398 213882 430634
rect 213326 394718 213562 394954
rect 213646 394718 213882 394954
rect 213326 394398 213562 394634
rect 213646 394398 213882 394634
rect 213326 358718 213562 358954
rect 213646 358718 213882 358954
rect 213326 358398 213562 358634
rect 213646 358398 213882 358634
rect 213326 322718 213562 322954
rect 213646 322718 213882 322954
rect 213326 322398 213562 322634
rect 213646 322398 213882 322634
rect 213326 286718 213562 286954
rect 213646 286718 213882 286954
rect 213326 286398 213562 286634
rect 213646 286398 213882 286634
rect 213326 250718 213562 250954
rect 213646 250718 213882 250954
rect 213326 250398 213562 250634
rect 213646 250398 213882 250634
rect 213326 214718 213562 214954
rect 213646 214718 213882 214954
rect 213326 214398 213562 214634
rect 213646 214398 213882 214634
rect 213326 178718 213562 178954
rect 213646 178718 213882 178954
rect 213326 178398 213562 178634
rect 213646 178398 213882 178634
rect 213326 142718 213562 142954
rect 213646 142718 213882 142954
rect 213326 142398 213562 142634
rect 213646 142398 213882 142634
rect 213326 106718 213562 106954
rect 213646 106718 213882 106954
rect 213326 106398 213562 106634
rect 213646 106398 213882 106634
rect 213326 70718 213562 70954
rect 213646 70718 213882 70954
rect 213326 70398 213562 70634
rect 213646 70398 213882 70634
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 222326 655718 222562 655954
rect 222646 655718 222882 655954
rect 222326 655398 222562 655634
rect 222646 655398 222882 655634
rect 222326 619718 222562 619954
rect 222646 619718 222882 619954
rect 222326 619398 222562 619634
rect 222646 619398 222882 619634
rect 222326 583718 222562 583954
rect 222646 583718 222882 583954
rect 222326 583398 222562 583634
rect 222646 583398 222882 583634
rect 222326 547718 222562 547954
rect 222646 547718 222882 547954
rect 222326 547398 222562 547634
rect 222646 547398 222882 547634
rect 222326 511718 222562 511954
rect 222646 511718 222882 511954
rect 222326 511398 222562 511634
rect 222646 511398 222882 511634
rect 222326 475718 222562 475954
rect 222646 475718 222882 475954
rect 222326 475398 222562 475634
rect 222646 475398 222882 475634
rect 222326 439718 222562 439954
rect 222646 439718 222882 439954
rect 222326 439398 222562 439634
rect 222646 439398 222882 439634
rect 222326 403718 222562 403954
rect 222646 403718 222882 403954
rect 222326 403398 222562 403634
rect 222646 403398 222882 403634
rect 222326 367718 222562 367954
rect 222646 367718 222882 367954
rect 222326 367398 222562 367634
rect 222646 367398 222882 367634
rect 222326 331718 222562 331954
rect 222646 331718 222882 331954
rect 222326 331398 222562 331634
rect 222646 331398 222882 331634
rect 222326 295718 222562 295954
rect 222646 295718 222882 295954
rect 222326 295398 222562 295634
rect 222646 295398 222882 295634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 222326 187718 222562 187954
rect 222646 187718 222882 187954
rect 222326 187398 222562 187634
rect 222646 187398 222882 187634
rect 222326 151718 222562 151954
rect 222646 151718 222882 151954
rect 222326 151398 222562 151634
rect 222646 151398 222882 151634
rect 222326 115718 222562 115954
rect 222646 115718 222882 115954
rect 222326 115398 222562 115634
rect 222646 115398 222882 115634
rect 222326 79718 222562 79954
rect 222646 79718 222882 79954
rect 222326 79398 222562 79634
rect 222646 79398 222882 79634
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 226826 660218 227062 660454
rect 227146 660218 227382 660454
rect 226826 659898 227062 660134
rect 227146 659898 227382 660134
rect 226826 624218 227062 624454
rect 227146 624218 227382 624454
rect 226826 623898 227062 624134
rect 227146 623898 227382 624134
rect 226826 588218 227062 588454
rect 227146 588218 227382 588454
rect 226826 587898 227062 588134
rect 227146 587898 227382 588134
rect 226826 552218 227062 552454
rect 227146 552218 227382 552454
rect 226826 551898 227062 552134
rect 227146 551898 227382 552134
rect 226826 516218 227062 516454
rect 227146 516218 227382 516454
rect 226826 515898 227062 516134
rect 227146 515898 227382 516134
rect 226826 480218 227062 480454
rect 227146 480218 227382 480454
rect 226826 479898 227062 480134
rect 227146 479898 227382 480134
rect 226826 444218 227062 444454
rect 227146 444218 227382 444454
rect 226826 443898 227062 444134
rect 227146 443898 227382 444134
rect 226826 408218 227062 408454
rect 227146 408218 227382 408454
rect 226826 407898 227062 408134
rect 227146 407898 227382 408134
rect 226826 372218 227062 372454
rect 227146 372218 227382 372454
rect 226826 371898 227062 372134
rect 227146 371898 227382 372134
rect 226826 336218 227062 336454
rect 227146 336218 227382 336454
rect 226826 335898 227062 336134
rect 227146 335898 227382 336134
rect 226826 300218 227062 300454
rect 227146 300218 227382 300454
rect 226826 299898 227062 300134
rect 227146 299898 227382 300134
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 231326 628718 231562 628954
rect 231646 628718 231882 628954
rect 231326 628398 231562 628634
rect 231646 628398 231882 628634
rect 231326 592718 231562 592954
rect 231646 592718 231882 592954
rect 231326 592398 231562 592634
rect 231646 592398 231882 592634
rect 231326 556718 231562 556954
rect 231646 556718 231882 556954
rect 231326 556398 231562 556634
rect 231646 556398 231882 556634
rect 231326 520718 231562 520954
rect 231646 520718 231882 520954
rect 231326 520398 231562 520634
rect 231646 520398 231882 520634
rect 231326 484718 231562 484954
rect 231646 484718 231882 484954
rect 231326 484398 231562 484634
rect 231646 484398 231882 484634
rect 231326 448718 231562 448954
rect 231646 448718 231882 448954
rect 231326 448398 231562 448634
rect 231646 448398 231882 448634
rect 231326 412718 231562 412954
rect 231646 412718 231882 412954
rect 231326 412398 231562 412634
rect 231646 412398 231882 412634
rect 231326 376718 231562 376954
rect 231646 376718 231882 376954
rect 231326 376398 231562 376634
rect 231646 376398 231882 376634
rect 231326 340718 231562 340954
rect 231646 340718 231882 340954
rect 231326 340398 231562 340634
rect 231646 340398 231882 340634
rect 231326 304718 231562 304954
rect 231646 304718 231882 304954
rect 231326 304398 231562 304634
rect 231646 304398 231882 304634
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 240326 637718 240562 637954
rect 240646 637718 240882 637954
rect 240326 637398 240562 637634
rect 240646 637398 240882 637634
rect 240326 601718 240562 601954
rect 240646 601718 240882 601954
rect 240326 601398 240562 601634
rect 240646 601398 240882 601634
rect 240326 565718 240562 565954
rect 240646 565718 240882 565954
rect 240326 565398 240562 565634
rect 240646 565398 240882 565634
rect 240326 529718 240562 529954
rect 240646 529718 240882 529954
rect 240326 529398 240562 529634
rect 240646 529398 240882 529634
rect 240326 493718 240562 493954
rect 240646 493718 240882 493954
rect 240326 493398 240562 493634
rect 240646 493398 240882 493634
rect 240326 457718 240562 457954
rect 240646 457718 240882 457954
rect 240326 457398 240562 457634
rect 240646 457398 240882 457634
rect 240326 421718 240562 421954
rect 240646 421718 240882 421954
rect 240326 421398 240562 421634
rect 240646 421398 240882 421634
rect 240326 385718 240562 385954
rect 240646 385718 240882 385954
rect 240326 385398 240562 385634
rect 240646 385398 240882 385634
rect 240326 349718 240562 349954
rect 240646 349718 240882 349954
rect 240326 349398 240562 349634
rect 240646 349398 240882 349634
rect 240326 313718 240562 313954
rect 240646 313718 240882 313954
rect 240326 313398 240562 313634
rect 240646 313398 240882 313634
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 244826 642218 245062 642454
rect 245146 642218 245382 642454
rect 244826 641898 245062 642134
rect 245146 641898 245382 642134
rect 244826 606218 245062 606454
rect 245146 606218 245382 606454
rect 244826 605898 245062 606134
rect 245146 605898 245382 606134
rect 244826 570218 245062 570454
rect 245146 570218 245382 570454
rect 244826 569898 245062 570134
rect 245146 569898 245382 570134
rect 244826 534218 245062 534454
rect 245146 534218 245382 534454
rect 244826 533898 245062 534134
rect 245146 533898 245382 534134
rect 244826 498218 245062 498454
rect 245146 498218 245382 498454
rect 244826 497898 245062 498134
rect 245146 497898 245382 498134
rect 244826 462218 245062 462454
rect 245146 462218 245382 462454
rect 244826 461898 245062 462134
rect 245146 461898 245382 462134
rect 244826 426218 245062 426454
rect 245146 426218 245382 426454
rect 244826 425898 245062 426134
rect 245146 425898 245382 426134
rect 244826 390218 245062 390454
rect 245146 390218 245382 390454
rect 244826 389898 245062 390134
rect 245146 389898 245382 390134
rect 244826 354218 245062 354454
rect 245146 354218 245382 354454
rect 244826 353898 245062 354134
rect 245146 353898 245382 354134
rect 244826 318218 245062 318454
rect 245146 318218 245382 318454
rect 244826 317898 245062 318134
rect 245146 317898 245382 318134
rect 244826 282218 245062 282454
rect 245146 282218 245382 282454
rect 244826 281898 245062 282134
rect 245146 281898 245382 282134
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 249326 646718 249562 646954
rect 249646 646718 249882 646954
rect 249326 646398 249562 646634
rect 249646 646398 249882 646634
rect 249326 610718 249562 610954
rect 249646 610718 249882 610954
rect 249326 610398 249562 610634
rect 249646 610398 249882 610634
rect 249326 574718 249562 574954
rect 249646 574718 249882 574954
rect 249326 574398 249562 574634
rect 249646 574398 249882 574634
rect 249326 538718 249562 538954
rect 249646 538718 249882 538954
rect 249326 538398 249562 538634
rect 249646 538398 249882 538634
rect 249326 502718 249562 502954
rect 249646 502718 249882 502954
rect 249326 502398 249562 502634
rect 249646 502398 249882 502634
rect 249326 466718 249562 466954
rect 249646 466718 249882 466954
rect 249326 466398 249562 466634
rect 249646 466398 249882 466634
rect 249326 430718 249562 430954
rect 249646 430718 249882 430954
rect 249326 430398 249562 430634
rect 249646 430398 249882 430634
rect 249326 394718 249562 394954
rect 249646 394718 249882 394954
rect 249326 394398 249562 394634
rect 249646 394398 249882 394634
rect 249326 358718 249562 358954
rect 249646 358718 249882 358954
rect 249326 358398 249562 358634
rect 249646 358398 249882 358634
rect 249326 322718 249562 322954
rect 249646 322718 249882 322954
rect 249326 322398 249562 322634
rect 249646 322398 249882 322634
rect 249326 286718 249562 286954
rect 249646 286718 249882 286954
rect 249326 286398 249562 286634
rect 249646 286398 249882 286634
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 276326 637718 276562 637954
rect 276646 637718 276882 637954
rect 276326 637398 276562 637634
rect 276646 637398 276882 637634
rect 276326 601718 276562 601954
rect 276646 601718 276882 601954
rect 276326 601398 276562 601634
rect 276646 601398 276882 601634
rect 276326 565718 276562 565954
rect 276646 565718 276882 565954
rect 276326 565398 276562 565634
rect 276646 565398 276882 565634
rect 276326 529718 276562 529954
rect 276646 529718 276882 529954
rect 276326 529398 276562 529634
rect 276646 529398 276882 529634
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 280826 642218 281062 642454
rect 281146 642218 281382 642454
rect 280826 641898 281062 642134
rect 281146 641898 281382 642134
rect 280826 606218 281062 606454
rect 281146 606218 281382 606454
rect 280826 605898 281062 606134
rect 281146 605898 281382 606134
rect 280826 570218 281062 570454
rect 281146 570218 281382 570454
rect 280826 569898 281062 570134
rect 281146 569898 281382 570134
rect 280826 534218 281062 534454
rect 281146 534218 281382 534454
rect 280826 533898 281062 534134
rect 281146 533898 281382 534134
rect 280826 498218 281062 498454
rect 281146 498218 281382 498454
rect 280826 497898 281062 498134
rect 281146 497898 281382 498134
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 285326 610718 285562 610954
rect 285646 610718 285882 610954
rect 285326 610398 285562 610634
rect 285646 610398 285882 610634
rect 285326 574718 285562 574954
rect 285646 574718 285882 574954
rect 285326 574398 285562 574634
rect 285646 574398 285882 574634
rect 285326 538718 285562 538954
rect 285646 538718 285882 538954
rect 285326 538398 285562 538634
rect 285646 538398 285882 538634
rect 285326 502718 285562 502954
rect 285646 502718 285882 502954
rect 285326 502398 285562 502634
rect 285646 502398 285882 502634
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 294326 619718 294562 619954
rect 294646 619718 294882 619954
rect 294326 619398 294562 619634
rect 294646 619398 294882 619634
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 294326 511718 294562 511954
rect 294646 511718 294882 511954
rect 294326 511398 294562 511634
rect 294646 511398 294882 511634
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 298826 624218 299062 624454
rect 299146 624218 299382 624454
rect 298826 623898 299062 624134
rect 299146 623898 299382 624134
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 298826 516218 299062 516454
rect 299146 516218 299382 516454
rect 298826 515898 299062 516134
rect 299146 515898 299382 516134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 298826 300218 299062 300454
rect 299146 300218 299382 300454
rect 298826 299898 299062 300134
rect 299146 299898 299382 300134
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 192218 299062 192454
rect 299146 192218 299382 192454
rect 298826 191898 299062 192134
rect 299146 191898 299382 192134
rect 298826 156218 299062 156454
rect 299146 156218 299382 156454
rect 298826 155898 299062 156134
rect 299146 155898 299382 156134
rect 298826 120218 299062 120454
rect 299146 120218 299382 120454
rect 298826 119898 299062 120134
rect 299146 119898 299382 120134
rect 298826 84218 299062 84454
rect 299146 84218 299382 84454
rect 298826 83898 299062 84134
rect 299146 83898 299382 84134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 303326 628718 303562 628954
rect 303646 628718 303882 628954
rect 303326 628398 303562 628634
rect 303646 628398 303882 628634
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 303326 520718 303562 520954
rect 303646 520718 303882 520954
rect 303326 520398 303562 520634
rect 303646 520398 303882 520634
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 303326 304718 303562 304954
rect 303646 304718 303882 304954
rect 303326 304398 303562 304634
rect 303646 304398 303882 304634
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 303326 196718 303562 196954
rect 303646 196718 303882 196954
rect 303326 196398 303562 196634
rect 303646 196398 303882 196634
rect 303326 160718 303562 160954
rect 303646 160718 303882 160954
rect 303326 160398 303562 160634
rect 303646 160398 303882 160634
rect 303326 124718 303562 124954
rect 303646 124718 303882 124954
rect 303326 124398 303562 124634
rect 303646 124398 303882 124634
rect 303326 88718 303562 88954
rect 303646 88718 303882 88954
rect 303326 88398 303562 88634
rect 303646 88398 303882 88634
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 312326 637718 312562 637954
rect 312646 637718 312882 637954
rect 312326 637398 312562 637634
rect 312646 637398 312882 637634
rect 312326 601718 312562 601954
rect 312646 601718 312882 601954
rect 312326 601398 312562 601634
rect 312646 601398 312882 601634
rect 312326 565718 312562 565954
rect 312646 565718 312882 565954
rect 312326 565398 312562 565634
rect 312646 565398 312882 565634
rect 312326 529718 312562 529954
rect 312646 529718 312882 529954
rect 312326 529398 312562 529634
rect 312646 529398 312882 529634
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 312326 313718 312562 313954
rect 312646 313718 312882 313954
rect 312326 313398 312562 313634
rect 312646 313398 312882 313634
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 312326 205718 312562 205954
rect 312646 205718 312882 205954
rect 312326 205398 312562 205634
rect 312646 205398 312882 205634
rect 312326 169718 312562 169954
rect 312646 169718 312882 169954
rect 312326 169398 312562 169634
rect 312646 169398 312882 169634
rect 312326 133718 312562 133954
rect 312646 133718 312882 133954
rect 312326 133398 312562 133634
rect 312646 133398 312882 133634
rect 312326 97718 312562 97954
rect 312646 97718 312882 97954
rect 312326 97398 312562 97634
rect 312646 97398 312882 97634
rect 312326 61718 312562 61954
rect 312646 61718 312882 61954
rect 312326 61398 312562 61634
rect 312646 61398 312882 61634
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 316826 642218 317062 642454
rect 317146 642218 317382 642454
rect 316826 641898 317062 642134
rect 317146 641898 317382 642134
rect 316826 606218 317062 606454
rect 317146 606218 317382 606454
rect 316826 605898 317062 606134
rect 317146 605898 317382 606134
rect 316826 570218 317062 570454
rect 317146 570218 317382 570454
rect 316826 569898 317062 570134
rect 317146 569898 317382 570134
rect 316826 534218 317062 534454
rect 317146 534218 317382 534454
rect 316826 533898 317062 534134
rect 317146 533898 317382 534134
rect 316826 498218 317062 498454
rect 317146 498218 317382 498454
rect 316826 497898 317062 498134
rect 317146 497898 317382 498134
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 316826 318218 317062 318454
rect 317146 318218 317382 318454
rect 316826 317898 317062 318134
rect 317146 317898 317382 318134
rect 316826 282218 317062 282454
rect 317146 282218 317382 282454
rect 316826 281898 317062 282134
rect 317146 281898 317382 282134
rect 316826 246218 317062 246454
rect 317146 246218 317382 246454
rect 316826 245898 317062 246134
rect 317146 245898 317382 246134
rect 316826 210218 317062 210454
rect 317146 210218 317382 210454
rect 316826 209898 317062 210134
rect 317146 209898 317382 210134
rect 316826 174218 317062 174454
rect 317146 174218 317382 174454
rect 316826 173898 317062 174134
rect 317146 173898 317382 174134
rect 316826 138218 317062 138454
rect 317146 138218 317382 138454
rect 316826 137898 317062 138134
rect 317146 137898 317382 138134
rect 316826 102218 317062 102454
rect 317146 102218 317382 102454
rect 316826 101898 317062 102134
rect 317146 101898 317382 102134
rect 316826 66218 317062 66454
rect 317146 66218 317382 66454
rect 316826 65898 317062 66134
rect 317146 65898 317382 66134
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 321326 610718 321562 610954
rect 321646 610718 321882 610954
rect 321326 610398 321562 610634
rect 321646 610398 321882 610634
rect 321326 574718 321562 574954
rect 321646 574718 321882 574954
rect 321326 574398 321562 574634
rect 321646 574398 321882 574634
rect 321326 538718 321562 538954
rect 321646 538718 321882 538954
rect 321326 538398 321562 538634
rect 321646 538398 321882 538634
rect 321326 502718 321562 502954
rect 321646 502718 321882 502954
rect 321326 502398 321562 502634
rect 321646 502398 321882 502634
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 321326 322718 321562 322954
rect 321646 322718 321882 322954
rect 321326 322398 321562 322634
rect 321646 322398 321882 322634
rect 321326 286718 321562 286954
rect 321646 286718 321882 286954
rect 321326 286398 321562 286634
rect 321646 286398 321882 286634
rect 321326 250718 321562 250954
rect 321646 250718 321882 250954
rect 321326 250398 321562 250634
rect 321646 250398 321882 250634
rect 321326 214718 321562 214954
rect 321646 214718 321882 214954
rect 321326 214398 321562 214634
rect 321646 214398 321882 214634
rect 321326 178718 321562 178954
rect 321646 178718 321882 178954
rect 321326 178398 321562 178634
rect 321646 178398 321882 178634
rect 321326 142718 321562 142954
rect 321646 142718 321882 142954
rect 321326 142398 321562 142634
rect 321646 142398 321882 142634
rect 321326 106718 321562 106954
rect 321646 106718 321882 106954
rect 321326 106398 321562 106634
rect 321646 106398 321882 106634
rect 321326 70718 321562 70954
rect 321646 70718 321882 70954
rect 321326 70398 321562 70634
rect 321646 70398 321882 70634
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 330326 331718 330562 331954
rect 330646 331718 330882 331954
rect 330326 331398 330562 331634
rect 330646 331398 330882 331634
rect 330326 295718 330562 295954
rect 330646 295718 330882 295954
rect 330326 295398 330562 295634
rect 330646 295398 330882 295634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 330326 187718 330562 187954
rect 330646 187718 330882 187954
rect 330326 187398 330562 187634
rect 330646 187398 330882 187634
rect 330326 151718 330562 151954
rect 330646 151718 330882 151954
rect 330326 151398 330562 151634
rect 330646 151398 330882 151634
rect 330326 115718 330562 115954
rect 330646 115718 330882 115954
rect 330326 115398 330562 115634
rect 330646 115398 330882 115634
rect 330326 79718 330562 79954
rect 330646 79718 330882 79954
rect 330326 79398 330562 79634
rect 330646 79398 330882 79634
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 334826 300218 335062 300454
rect 335146 300218 335382 300454
rect 334826 299898 335062 300134
rect 335146 299898 335382 300134
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 334826 192218 335062 192454
rect 335146 192218 335382 192454
rect 334826 191898 335062 192134
rect 335146 191898 335382 192134
rect 334826 156218 335062 156454
rect 335146 156218 335382 156454
rect 334826 155898 335062 156134
rect 335146 155898 335382 156134
rect 334826 120218 335062 120454
rect 335146 120218 335382 120454
rect 334826 119898 335062 120134
rect 335146 119898 335382 120134
rect 334826 84218 335062 84454
rect 335146 84218 335382 84454
rect 334826 83898 335062 84134
rect 335146 83898 335382 84134
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 339326 304718 339562 304954
rect 339646 304718 339882 304954
rect 339326 304398 339562 304634
rect 339646 304398 339882 304634
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 339326 196718 339562 196954
rect 339646 196718 339882 196954
rect 339326 196398 339562 196634
rect 339646 196398 339882 196634
rect 339326 160718 339562 160954
rect 339646 160718 339882 160954
rect 339326 160398 339562 160634
rect 339646 160398 339882 160634
rect 339326 124718 339562 124954
rect 339646 124718 339882 124954
rect 339326 124398 339562 124634
rect 339646 124398 339882 124634
rect 339326 88718 339562 88954
rect 339646 88718 339882 88954
rect 339326 88398 339562 88634
rect 339646 88398 339882 88634
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 348326 313718 348562 313954
rect 348646 313718 348882 313954
rect 348326 313398 348562 313634
rect 348646 313398 348882 313634
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 318218 353062 318454
rect 353146 318218 353382 318454
rect 352826 317898 353062 318134
rect 353146 317898 353382 318134
rect 352826 282218 353062 282454
rect 353146 282218 353382 282454
rect 352826 281898 353062 282134
rect 353146 281898 353382 282134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 357326 610718 357562 610954
rect 357646 610718 357882 610954
rect 357326 610398 357562 610634
rect 357646 610398 357882 610634
rect 357326 574718 357562 574954
rect 357646 574718 357882 574954
rect 357326 574398 357562 574634
rect 357646 574398 357882 574634
rect 357326 538718 357562 538954
rect 357646 538718 357882 538954
rect 357326 538398 357562 538634
rect 357646 538398 357882 538634
rect 357326 502718 357562 502954
rect 357646 502718 357882 502954
rect 357326 502398 357562 502634
rect 357646 502398 357882 502634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 366326 619718 366562 619954
rect 366646 619718 366882 619954
rect 366326 619398 366562 619634
rect 366646 619398 366882 619634
rect 366326 583718 366562 583954
rect 366646 583718 366882 583954
rect 366326 583398 366562 583634
rect 366646 583398 366882 583634
rect 366326 547718 366562 547954
rect 366646 547718 366882 547954
rect 366326 547398 366562 547634
rect 366646 547398 366882 547634
rect 366326 511718 366562 511954
rect 366646 511718 366882 511954
rect 366326 511398 366562 511634
rect 366646 511398 366882 511634
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 370826 624218 371062 624454
rect 371146 624218 371382 624454
rect 370826 623898 371062 624134
rect 371146 623898 371382 624134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 370826 552218 371062 552454
rect 371146 552218 371382 552454
rect 370826 551898 371062 552134
rect 371146 551898 371382 552134
rect 370826 516218 371062 516454
rect 371146 516218 371382 516454
rect 370826 515898 371062 516134
rect 371146 515898 371382 516134
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 375326 628718 375562 628954
rect 375646 628718 375882 628954
rect 375326 628398 375562 628634
rect 375646 628398 375882 628634
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 375326 520718 375562 520954
rect 375646 520718 375882 520954
rect 375326 520398 375562 520634
rect 375646 520398 375882 520634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 384326 637718 384562 637954
rect 384646 637718 384882 637954
rect 384326 637398 384562 637634
rect 384646 637398 384882 637634
rect 384326 601718 384562 601954
rect 384646 601718 384882 601954
rect 384326 601398 384562 601634
rect 384646 601398 384882 601634
rect 384326 565718 384562 565954
rect 384646 565718 384882 565954
rect 384326 565398 384562 565634
rect 384646 565398 384882 565634
rect 384326 529718 384562 529954
rect 384646 529718 384882 529954
rect 384326 529398 384562 529634
rect 384646 529398 384882 529634
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642218 389062 642454
rect 389146 642218 389382 642454
rect 388826 641898 389062 642134
rect 389146 641898 389382 642134
rect 388826 606218 389062 606454
rect 389146 606218 389382 606454
rect 388826 605898 389062 606134
rect 389146 605898 389382 606134
rect 388826 570218 389062 570454
rect 389146 570218 389382 570454
rect 388826 569898 389062 570134
rect 389146 569898 389382 570134
rect 388826 534218 389062 534454
rect 389146 534218 389382 534454
rect 388826 533898 389062 534134
rect 389146 533898 389382 534134
rect 388826 498218 389062 498454
rect 389146 498218 389382 498454
rect 388826 497898 389062 498134
rect 389146 497898 389382 498134
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 393326 610718 393562 610954
rect 393646 610718 393882 610954
rect 393326 610398 393562 610634
rect 393646 610398 393882 610634
rect 393326 574718 393562 574954
rect 393646 574718 393882 574954
rect 393326 574398 393562 574634
rect 393646 574398 393882 574634
rect 393326 538718 393562 538954
rect 393646 538718 393882 538954
rect 393326 538398 393562 538634
rect 393646 538398 393882 538634
rect 393326 502718 393562 502954
rect 393646 502718 393882 502954
rect 393326 502398 393562 502634
rect 393646 502398 393882 502634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 402326 619718 402562 619954
rect 402646 619718 402882 619954
rect 402326 619398 402562 619634
rect 402646 619398 402882 619634
rect 402326 583718 402562 583954
rect 402646 583718 402882 583954
rect 402326 583398 402562 583634
rect 402646 583398 402882 583634
rect 402326 547718 402562 547954
rect 402646 547718 402882 547954
rect 402326 547398 402562 547634
rect 402646 547398 402882 547634
rect 402326 511718 402562 511954
rect 402646 511718 402882 511954
rect 402326 511398 402562 511634
rect 402646 511398 402882 511634
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 478826 624218 479062 624454
rect 479146 624218 479382 624454
rect 478826 623898 479062 624134
rect 479146 623898 479382 624134
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 478826 516218 479062 516454
rect 479146 516218 479382 516454
rect 478826 515898 479062 516134
rect 479146 515898 479382 516134
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 483326 628718 483562 628954
rect 483646 628718 483882 628954
rect 483326 628398 483562 628634
rect 483646 628398 483882 628634
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 483326 520718 483562 520954
rect 483646 520718 483882 520954
rect 483326 520398 483562 520634
rect 483646 520398 483882 520634
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 492326 637718 492562 637954
rect 492646 637718 492882 637954
rect 492326 637398 492562 637634
rect 492646 637398 492882 637634
rect 492326 601718 492562 601954
rect 492646 601718 492882 601954
rect 492326 601398 492562 601634
rect 492646 601398 492882 601634
rect 492326 565718 492562 565954
rect 492646 565718 492882 565954
rect 492326 565398 492562 565634
rect 492646 565398 492882 565634
rect 492326 529718 492562 529954
rect 492646 529718 492882 529954
rect 492326 529398 492562 529634
rect 492646 529398 492882 529634
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642218 497062 642454
rect 497146 642218 497382 642454
rect 496826 641898 497062 642134
rect 497146 641898 497382 642134
rect 496826 606218 497062 606454
rect 497146 606218 497382 606454
rect 496826 605898 497062 606134
rect 497146 605898 497382 606134
rect 496826 570218 497062 570454
rect 497146 570218 497382 570454
rect 496826 569898 497062 570134
rect 497146 569898 497382 570134
rect 496826 534218 497062 534454
rect 497146 534218 497382 534454
rect 496826 533898 497062 534134
rect 497146 533898 497382 534134
rect 496826 498218 497062 498454
rect 497146 498218 497382 498454
rect 496826 497898 497062 498134
rect 497146 497898 497382 498134
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 501326 610718 501562 610954
rect 501646 610718 501882 610954
rect 501326 610398 501562 610634
rect 501646 610398 501882 610634
rect 501326 574718 501562 574954
rect 501646 574718 501882 574954
rect 501326 574398 501562 574634
rect 501646 574398 501882 574634
rect 501326 538718 501562 538954
rect 501646 538718 501882 538954
rect 501326 538398 501562 538634
rect 501646 538398 501882 538634
rect 501326 502718 501562 502954
rect 501646 502718 501882 502954
rect 501326 502398 501562 502634
rect 501646 502398 501882 502634
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 510326 619718 510562 619954
rect 510646 619718 510882 619954
rect 510326 619398 510562 619634
rect 510646 619398 510882 619634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 510326 511718 510562 511954
rect 510646 511718 510882 511954
rect 510326 511398 510562 511634
rect 510646 511398 510882 511634
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 514826 624218 515062 624454
rect 515146 624218 515382 624454
rect 514826 623898 515062 624134
rect 515146 623898 515382 624134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 514826 516218 515062 516454
rect 515146 516218 515382 516454
rect 514826 515898 515062 516134
rect 515146 515898 515382 516134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 519326 628718 519562 628954
rect 519646 628718 519882 628954
rect 519326 628398 519562 628634
rect 519646 628398 519882 628634
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 519326 520718 519562 520954
rect 519646 520718 519882 520954
rect 519326 520398 519562 520634
rect 519646 520398 519882 520634
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 82826 660454
rect 83062 660218 83146 660454
rect 83382 660218 118826 660454
rect 119062 660218 119146 660454
rect 119382 660218 154826 660454
rect 155062 660218 155146 660454
rect 155382 660218 190826 660454
rect 191062 660218 191146 660454
rect 191382 660218 226826 660454
rect 227062 660218 227146 660454
rect 227382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 82826 660134
rect 83062 659898 83146 660134
rect 83382 659898 118826 660134
rect 119062 659898 119146 660134
rect 119382 659898 154826 660134
rect 155062 659898 155146 660134
rect 155382 659898 190826 660134
rect 191062 659898 191146 660134
rect 191382 659898 226826 660134
rect 227062 659898 227146 660134
rect 227382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 78326 655954
rect 78562 655718 78646 655954
rect 78882 655718 114326 655954
rect 114562 655718 114646 655954
rect 114882 655718 150326 655954
rect 150562 655718 150646 655954
rect 150882 655718 186326 655954
rect 186562 655718 186646 655954
rect 186882 655718 222326 655954
rect 222562 655718 222646 655954
rect 222882 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 78326 655634
rect 78562 655398 78646 655634
rect 78882 655398 114326 655634
rect 114562 655398 114646 655634
rect 114882 655398 150326 655634
rect 150562 655398 150646 655634
rect 150882 655398 186326 655634
rect 186562 655398 186646 655634
rect 186882 655398 222326 655634
rect 222562 655398 222646 655634
rect 222882 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 69326 646954
rect 69562 646718 69646 646954
rect 69882 646718 105326 646954
rect 105562 646718 105646 646954
rect 105882 646718 141326 646954
rect 141562 646718 141646 646954
rect 141882 646718 177326 646954
rect 177562 646718 177646 646954
rect 177882 646718 213326 646954
rect 213562 646718 213646 646954
rect 213882 646718 249326 646954
rect 249562 646718 249646 646954
rect 249882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 69326 646634
rect 69562 646398 69646 646634
rect 69882 646398 105326 646634
rect 105562 646398 105646 646634
rect 105882 646398 141326 646634
rect 141562 646398 141646 646634
rect 141882 646398 177326 646634
rect 177562 646398 177646 646634
rect 177882 646398 213326 646634
rect 213562 646398 213646 646634
rect 213882 646398 249326 646634
rect 249562 646398 249646 646634
rect 249882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 64826 642454
rect 65062 642218 65146 642454
rect 65382 642218 100826 642454
rect 101062 642218 101146 642454
rect 101382 642218 136826 642454
rect 137062 642218 137146 642454
rect 137382 642218 172826 642454
rect 173062 642218 173146 642454
rect 173382 642218 208826 642454
rect 209062 642218 209146 642454
rect 209382 642218 244826 642454
rect 245062 642218 245146 642454
rect 245382 642218 280826 642454
rect 281062 642218 281146 642454
rect 281382 642218 316826 642454
rect 317062 642218 317146 642454
rect 317382 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 388826 642454
rect 389062 642218 389146 642454
rect 389382 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 496826 642454
rect 497062 642218 497146 642454
rect 497382 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect -8726 642134 592650 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 64826 642134
rect 65062 641898 65146 642134
rect 65382 641898 100826 642134
rect 101062 641898 101146 642134
rect 101382 641898 136826 642134
rect 137062 641898 137146 642134
rect 137382 641898 172826 642134
rect 173062 641898 173146 642134
rect 173382 641898 208826 642134
rect 209062 641898 209146 642134
rect 209382 641898 244826 642134
rect 245062 641898 245146 642134
rect 245382 641898 280826 642134
rect 281062 641898 281146 642134
rect 281382 641898 316826 642134
rect 317062 641898 317146 642134
rect 317382 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 388826 642134
rect 389062 641898 389146 642134
rect 389382 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 496826 642134
rect 497062 641898 497146 642134
rect 497382 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 60326 637954
rect 60562 637718 60646 637954
rect 60882 637718 96326 637954
rect 96562 637718 96646 637954
rect 96882 637718 132326 637954
rect 132562 637718 132646 637954
rect 132882 637718 168326 637954
rect 168562 637718 168646 637954
rect 168882 637718 204326 637954
rect 204562 637718 204646 637954
rect 204882 637718 240326 637954
rect 240562 637718 240646 637954
rect 240882 637718 276326 637954
rect 276562 637718 276646 637954
rect 276882 637718 312326 637954
rect 312562 637718 312646 637954
rect 312882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 384326 637954
rect 384562 637718 384646 637954
rect 384882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 492326 637954
rect 492562 637718 492646 637954
rect 492882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 60326 637634
rect 60562 637398 60646 637634
rect 60882 637398 96326 637634
rect 96562 637398 96646 637634
rect 96882 637398 132326 637634
rect 132562 637398 132646 637634
rect 132882 637398 168326 637634
rect 168562 637398 168646 637634
rect 168882 637398 204326 637634
rect 204562 637398 204646 637634
rect 204882 637398 240326 637634
rect 240562 637398 240646 637634
rect 240882 637398 276326 637634
rect 276562 637398 276646 637634
rect 276882 637398 312326 637634
rect 312562 637398 312646 637634
rect 312882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 384326 637634
rect 384562 637398 384646 637634
rect 384882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 492326 637634
rect 492562 637398 492646 637634
rect 492882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 51326 628954
rect 51562 628718 51646 628954
rect 51882 628718 87326 628954
rect 87562 628718 87646 628954
rect 87882 628718 123326 628954
rect 123562 628718 123646 628954
rect 123882 628718 159326 628954
rect 159562 628718 159646 628954
rect 159882 628718 195326 628954
rect 195562 628718 195646 628954
rect 195882 628718 231326 628954
rect 231562 628718 231646 628954
rect 231882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 303326 628954
rect 303562 628718 303646 628954
rect 303882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 375326 628954
rect 375562 628718 375646 628954
rect 375882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 483326 628954
rect 483562 628718 483646 628954
rect 483882 628718 519326 628954
rect 519562 628718 519646 628954
rect 519882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 51326 628634
rect 51562 628398 51646 628634
rect 51882 628398 87326 628634
rect 87562 628398 87646 628634
rect 87882 628398 123326 628634
rect 123562 628398 123646 628634
rect 123882 628398 159326 628634
rect 159562 628398 159646 628634
rect 159882 628398 195326 628634
rect 195562 628398 195646 628634
rect 195882 628398 231326 628634
rect 231562 628398 231646 628634
rect 231882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 303326 628634
rect 303562 628398 303646 628634
rect 303882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 375326 628634
rect 375562 628398 375646 628634
rect 375882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 483326 628634
rect 483562 628398 483646 628634
rect 483882 628398 519326 628634
rect 519562 628398 519646 628634
rect 519882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 82826 624454
rect 83062 624218 83146 624454
rect 83382 624218 118826 624454
rect 119062 624218 119146 624454
rect 119382 624218 154826 624454
rect 155062 624218 155146 624454
rect 155382 624218 190826 624454
rect 191062 624218 191146 624454
rect 191382 624218 226826 624454
rect 227062 624218 227146 624454
rect 227382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 298826 624454
rect 299062 624218 299146 624454
rect 299382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 370826 624454
rect 371062 624218 371146 624454
rect 371382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 478826 624454
rect 479062 624218 479146 624454
rect 479382 624218 514826 624454
rect 515062 624218 515146 624454
rect 515382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 82826 624134
rect 83062 623898 83146 624134
rect 83382 623898 118826 624134
rect 119062 623898 119146 624134
rect 119382 623898 154826 624134
rect 155062 623898 155146 624134
rect 155382 623898 190826 624134
rect 191062 623898 191146 624134
rect 191382 623898 226826 624134
rect 227062 623898 227146 624134
rect 227382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 298826 624134
rect 299062 623898 299146 624134
rect 299382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 370826 624134
rect 371062 623898 371146 624134
rect 371382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 478826 624134
rect 479062 623898 479146 624134
rect 479382 623898 514826 624134
rect 515062 623898 515146 624134
rect 515382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 78326 619954
rect 78562 619718 78646 619954
rect 78882 619718 114326 619954
rect 114562 619718 114646 619954
rect 114882 619718 150326 619954
rect 150562 619718 150646 619954
rect 150882 619718 186326 619954
rect 186562 619718 186646 619954
rect 186882 619718 222326 619954
rect 222562 619718 222646 619954
rect 222882 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 294326 619954
rect 294562 619718 294646 619954
rect 294882 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 366326 619954
rect 366562 619718 366646 619954
rect 366882 619718 402326 619954
rect 402562 619718 402646 619954
rect 402882 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 510326 619954
rect 510562 619718 510646 619954
rect 510882 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 78326 619634
rect 78562 619398 78646 619634
rect 78882 619398 114326 619634
rect 114562 619398 114646 619634
rect 114882 619398 150326 619634
rect 150562 619398 150646 619634
rect 150882 619398 186326 619634
rect 186562 619398 186646 619634
rect 186882 619398 222326 619634
rect 222562 619398 222646 619634
rect 222882 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 294326 619634
rect 294562 619398 294646 619634
rect 294882 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 366326 619634
rect 366562 619398 366646 619634
rect 366882 619398 402326 619634
rect 402562 619398 402646 619634
rect 402882 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 510326 619634
rect 510562 619398 510646 619634
rect 510882 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 69326 610954
rect 69562 610718 69646 610954
rect 69882 610718 105326 610954
rect 105562 610718 105646 610954
rect 105882 610718 141326 610954
rect 141562 610718 141646 610954
rect 141882 610718 177326 610954
rect 177562 610718 177646 610954
rect 177882 610718 213326 610954
rect 213562 610718 213646 610954
rect 213882 610718 249326 610954
rect 249562 610718 249646 610954
rect 249882 610718 285326 610954
rect 285562 610718 285646 610954
rect 285882 610718 321326 610954
rect 321562 610718 321646 610954
rect 321882 610718 357326 610954
rect 357562 610718 357646 610954
rect 357882 610718 393326 610954
rect 393562 610718 393646 610954
rect 393882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 501326 610954
rect 501562 610718 501646 610954
rect 501882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 69326 610634
rect 69562 610398 69646 610634
rect 69882 610398 105326 610634
rect 105562 610398 105646 610634
rect 105882 610398 141326 610634
rect 141562 610398 141646 610634
rect 141882 610398 177326 610634
rect 177562 610398 177646 610634
rect 177882 610398 213326 610634
rect 213562 610398 213646 610634
rect 213882 610398 249326 610634
rect 249562 610398 249646 610634
rect 249882 610398 285326 610634
rect 285562 610398 285646 610634
rect 285882 610398 321326 610634
rect 321562 610398 321646 610634
rect 321882 610398 357326 610634
rect 357562 610398 357646 610634
rect 357882 610398 393326 610634
rect 393562 610398 393646 610634
rect 393882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 501326 610634
rect 501562 610398 501646 610634
rect 501882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 64826 606454
rect 65062 606218 65146 606454
rect 65382 606218 100826 606454
rect 101062 606218 101146 606454
rect 101382 606218 136826 606454
rect 137062 606218 137146 606454
rect 137382 606218 172826 606454
rect 173062 606218 173146 606454
rect 173382 606218 208826 606454
rect 209062 606218 209146 606454
rect 209382 606218 244826 606454
rect 245062 606218 245146 606454
rect 245382 606218 280826 606454
rect 281062 606218 281146 606454
rect 281382 606218 316826 606454
rect 317062 606218 317146 606454
rect 317382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 388826 606454
rect 389062 606218 389146 606454
rect 389382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 496826 606454
rect 497062 606218 497146 606454
rect 497382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 64826 606134
rect 65062 605898 65146 606134
rect 65382 605898 100826 606134
rect 101062 605898 101146 606134
rect 101382 605898 136826 606134
rect 137062 605898 137146 606134
rect 137382 605898 172826 606134
rect 173062 605898 173146 606134
rect 173382 605898 208826 606134
rect 209062 605898 209146 606134
rect 209382 605898 244826 606134
rect 245062 605898 245146 606134
rect 245382 605898 280826 606134
rect 281062 605898 281146 606134
rect 281382 605898 316826 606134
rect 317062 605898 317146 606134
rect 317382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 388826 606134
rect 389062 605898 389146 606134
rect 389382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 496826 606134
rect 497062 605898 497146 606134
rect 497382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 60326 601954
rect 60562 601718 60646 601954
rect 60882 601718 96326 601954
rect 96562 601718 96646 601954
rect 96882 601718 132326 601954
rect 132562 601718 132646 601954
rect 132882 601718 168326 601954
rect 168562 601718 168646 601954
rect 168882 601718 204326 601954
rect 204562 601718 204646 601954
rect 204882 601718 240326 601954
rect 240562 601718 240646 601954
rect 240882 601718 276326 601954
rect 276562 601718 276646 601954
rect 276882 601718 312326 601954
rect 312562 601718 312646 601954
rect 312882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 384326 601954
rect 384562 601718 384646 601954
rect 384882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 492326 601954
rect 492562 601718 492646 601954
rect 492882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 60326 601634
rect 60562 601398 60646 601634
rect 60882 601398 96326 601634
rect 96562 601398 96646 601634
rect 96882 601398 132326 601634
rect 132562 601398 132646 601634
rect 132882 601398 168326 601634
rect 168562 601398 168646 601634
rect 168882 601398 204326 601634
rect 204562 601398 204646 601634
rect 204882 601398 240326 601634
rect 240562 601398 240646 601634
rect 240882 601398 276326 601634
rect 276562 601398 276646 601634
rect 276882 601398 312326 601634
rect 312562 601398 312646 601634
rect 312882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 384326 601634
rect 384562 601398 384646 601634
rect 384882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 492326 601634
rect 492562 601398 492646 601634
rect 492882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 51326 592954
rect 51562 592718 51646 592954
rect 51882 592718 87326 592954
rect 87562 592718 87646 592954
rect 87882 592718 123326 592954
rect 123562 592718 123646 592954
rect 123882 592718 159326 592954
rect 159562 592718 159646 592954
rect 159882 592718 195326 592954
rect 195562 592718 195646 592954
rect 195882 592718 231326 592954
rect 231562 592718 231646 592954
rect 231882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 51326 592634
rect 51562 592398 51646 592634
rect 51882 592398 87326 592634
rect 87562 592398 87646 592634
rect 87882 592398 123326 592634
rect 123562 592398 123646 592634
rect 123882 592398 159326 592634
rect 159562 592398 159646 592634
rect 159882 592398 195326 592634
rect 195562 592398 195646 592634
rect 195882 592398 231326 592634
rect 231562 592398 231646 592634
rect 231882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 82826 588454
rect 83062 588218 83146 588454
rect 83382 588218 118826 588454
rect 119062 588218 119146 588454
rect 119382 588218 154826 588454
rect 155062 588218 155146 588454
rect 155382 588218 190826 588454
rect 191062 588218 191146 588454
rect 191382 588218 226826 588454
rect 227062 588218 227146 588454
rect 227382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 82826 588134
rect 83062 587898 83146 588134
rect 83382 587898 118826 588134
rect 119062 587898 119146 588134
rect 119382 587898 154826 588134
rect 155062 587898 155146 588134
rect 155382 587898 190826 588134
rect 191062 587898 191146 588134
rect 191382 587898 226826 588134
rect 227062 587898 227146 588134
rect 227382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 78326 583954
rect 78562 583718 78646 583954
rect 78882 583718 114326 583954
rect 114562 583718 114646 583954
rect 114882 583718 150326 583954
rect 150562 583718 150646 583954
rect 150882 583718 186326 583954
rect 186562 583718 186646 583954
rect 186882 583718 222326 583954
rect 222562 583718 222646 583954
rect 222882 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 366326 583954
rect 366562 583718 366646 583954
rect 366882 583718 402326 583954
rect 402562 583718 402646 583954
rect 402882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 78326 583634
rect 78562 583398 78646 583634
rect 78882 583398 114326 583634
rect 114562 583398 114646 583634
rect 114882 583398 150326 583634
rect 150562 583398 150646 583634
rect 150882 583398 186326 583634
rect 186562 583398 186646 583634
rect 186882 583398 222326 583634
rect 222562 583398 222646 583634
rect 222882 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 366326 583634
rect 366562 583398 366646 583634
rect 366882 583398 402326 583634
rect 402562 583398 402646 583634
rect 402882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 69326 574954
rect 69562 574718 69646 574954
rect 69882 574718 105326 574954
rect 105562 574718 105646 574954
rect 105882 574718 141326 574954
rect 141562 574718 141646 574954
rect 141882 574718 177326 574954
rect 177562 574718 177646 574954
rect 177882 574718 213326 574954
rect 213562 574718 213646 574954
rect 213882 574718 249326 574954
rect 249562 574718 249646 574954
rect 249882 574718 285326 574954
rect 285562 574718 285646 574954
rect 285882 574718 321326 574954
rect 321562 574718 321646 574954
rect 321882 574718 357326 574954
rect 357562 574718 357646 574954
rect 357882 574718 393326 574954
rect 393562 574718 393646 574954
rect 393882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 501326 574954
rect 501562 574718 501646 574954
rect 501882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 69326 574634
rect 69562 574398 69646 574634
rect 69882 574398 105326 574634
rect 105562 574398 105646 574634
rect 105882 574398 141326 574634
rect 141562 574398 141646 574634
rect 141882 574398 177326 574634
rect 177562 574398 177646 574634
rect 177882 574398 213326 574634
rect 213562 574398 213646 574634
rect 213882 574398 249326 574634
rect 249562 574398 249646 574634
rect 249882 574398 285326 574634
rect 285562 574398 285646 574634
rect 285882 574398 321326 574634
rect 321562 574398 321646 574634
rect 321882 574398 357326 574634
rect 357562 574398 357646 574634
rect 357882 574398 393326 574634
rect 393562 574398 393646 574634
rect 393882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 501326 574634
rect 501562 574398 501646 574634
rect 501882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 64826 570454
rect 65062 570218 65146 570454
rect 65382 570218 100826 570454
rect 101062 570218 101146 570454
rect 101382 570218 136826 570454
rect 137062 570218 137146 570454
rect 137382 570218 172826 570454
rect 173062 570218 173146 570454
rect 173382 570218 208826 570454
rect 209062 570218 209146 570454
rect 209382 570218 244826 570454
rect 245062 570218 245146 570454
rect 245382 570218 280826 570454
rect 281062 570218 281146 570454
rect 281382 570218 316826 570454
rect 317062 570218 317146 570454
rect 317382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 388826 570454
rect 389062 570218 389146 570454
rect 389382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 496826 570454
rect 497062 570218 497146 570454
rect 497382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 64826 570134
rect 65062 569898 65146 570134
rect 65382 569898 100826 570134
rect 101062 569898 101146 570134
rect 101382 569898 136826 570134
rect 137062 569898 137146 570134
rect 137382 569898 172826 570134
rect 173062 569898 173146 570134
rect 173382 569898 208826 570134
rect 209062 569898 209146 570134
rect 209382 569898 244826 570134
rect 245062 569898 245146 570134
rect 245382 569898 280826 570134
rect 281062 569898 281146 570134
rect 281382 569898 316826 570134
rect 317062 569898 317146 570134
rect 317382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 388826 570134
rect 389062 569898 389146 570134
rect 389382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 496826 570134
rect 497062 569898 497146 570134
rect 497382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 60326 565954
rect 60562 565718 60646 565954
rect 60882 565718 96326 565954
rect 96562 565718 96646 565954
rect 96882 565718 132326 565954
rect 132562 565718 132646 565954
rect 132882 565718 168326 565954
rect 168562 565718 168646 565954
rect 168882 565718 204326 565954
rect 204562 565718 204646 565954
rect 204882 565718 240326 565954
rect 240562 565718 240646 565954
rect 240882 565718 276326 565954
rect 276562 565718 276646 565954
rect 276882 565718 312326 565954
rect 312562 565718 312646 565954
rect 312882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 384326 565954
rect 384562 565718 384646 565954
rect 384882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 492326 565954
rect 492562 565718 492646 565954
rect 492882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 60326 565634
rect 60562 565398 60646 565634
rect 60882 565398 96326 565634
rect 96562 565398 96646 565634
rect 96882 565398 132326 565634
rect 132562 565398 132646 565634
rect 132882 565398 168326 565634
rect 168562 565398 168646 565634
rect 168882 565398 204326 565634
rect 204562 565398 204646 565634
rect 204882 565398 240326 565634
rect 240562 565398 240646 565634
rect 240882 565398 276326 565634
rect 276562 565398 276646 565634
rect 276882 565398 312326 565634
rect 312562 565398 312646 565634
rect 312882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 384326 565634
rect 384562 565398 384646 565634
rect 384882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 492326 565634
rect 492562 565398 492646 565634
rect 492882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 51326 556954
rect 51562 556718 51646 556954
rect 51882 556718 87326 556954
rect 87562 556718 87646 556954
rect 87882 556718 123326 556954
rect 123562 556718 123646 556954
rect 123882 556718 159326 556954
rect 159562 556718 159646 556954
rect 159882 556718 195326 556954
rect 195562 556718 195646 556954
rect 195882 556718 231326 556954
rect 231562 556718 231646 556954
rect 231882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 51326 556634
rect 51562 556398 51646 556634
rect 51882 556398 87326 556634
rect 87562 556398 87646 556634
rect 87882 556398 123326 556634
rect 123562 556398 123646 556634
rect 123882 556398 159326 556634
rect 159562 556398 159646 556634
rect 159882 556398 195326 556634
rect 195562 556398 195646 556634
rect 195882 556398 231326 556634
rect 231562 556398 231646 556634
rect 231882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 82826 552454
rect 83062 552218 83146 552454
rect 83382 552218 118826 552454
rect 119062 552218 119146 552454
rect 119382 552218 154826 552454
rect 155062 552218 155146 552454
rect 155382 552218 190826 552454
rect 191062 552218 191146 552454
rect 191382 552218 226826 552454
rect 227062 552218 227146 552454
rect 227382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 370826 552454
rect 371062 552218 371146 552454
rect 371382 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 82826 552134
rect 83062 551898 83146 552134
rect 83382 551898 118826 552134
rect 119062 551898 119146 552134
rect 119382 551898 154826 552134
rect 155062 551898 155146 552134
rect 155382 551898 190826 552134
rect 191062 551898 191146 552134
rect 191382 551898 226826 552134
rect 227062 551898 227146 552134
rect 227382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 370826 552134
rect 371062 551898 371146 552134
rect 371382 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 78326 547954
rect 78562 547718 78646 547954
rect 78882 547718 114326 547954
rect 114562 547718 114646 547954
rect 114882 547718 150326 547954
rect 150562 547718 150646 547954
rect 150882 547718 186326 547954
rect 186562 547718 186646 547954
rect 186882 547718 222326 547954
rect 222562 547718 222646 547954
rect 222882 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 366326 547954
rect 366562 547718 366646 547954
rect 366882 547718 402326 547954
rect 402562 547718 402646 547954
rect 402882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 78326 547634
rect 78562 547398 78646 547634
rect 78882 547398 114326 547634
rect 114562 547398 114646 547634
rect 114882 547398 150326 547634
rect 150562 547398 150646 547634
rect 150882 547398 186326 547634
rect 186562 547398 186646 547634
rect 186882 547398 222326 547634
rect 222562 547398 222646 547634
rect 222882 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 366326 547634
rect 366562 547398 366646 547634
rect 366882 547398 402326 547634
rect 402562 547398 402646 547634
rect 402882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 69326 538954
rect 69562 538718 69646 538954
rect 69882 538718 105326 538954
rect 105562 538718 105646 538954
rect 105882 538718 141326 538954
rect 141562 538718 141646 538954
rect 141882 538718 177326 538954
rect 177562 538718 177646 538954
rect 177882 538718 213326 538954
rect 213562 538718 213646 538954
rect 213882 538718 249326 538954
rect 249562 538718 249646 538954
rect 249882 538718 285326 538954
rect 285562 538718 285646 538954
rect 285882 538718 321326 538954
rect 321562 538718 321646 538954
rect 321882 538718 357326 538954
rect 357562 538718 357646 538954
rect 357882 538718 393326 538954
rect 393562 538718 393646 538954
rect 393882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 501326 538954
rect 501562 538718 501646 538954
rect 501882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 69326 538634
rect 69562 538398 69646 538634
rect 69882 538398 105326 538634
rect 105562 538398 105646 538634
rect 105882 538398 141326 538634
rect 141562 538398 141646 538634
rect 141882 538398 177326 538634
rect 177562 538398 177646 538634
rect 177882 538398 213326 538634
rect 213562 538398 213646 538634
rect 213882 538398 249326 538634
rect 249562 538398 249646 538634
rect 249882 538398 285326 538634
rect 285562 538398 285646 538634
rect 285882 538398 321326 538634
rect 321562 538398 321646 538634
rect 321882 538398 357326 538634
rect 357562 538398 357646 538634
rect 357882 538398 393326 538634
rect 393562 538398 393646 538634
rect 393882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 501326 538634
rect 501562 538398 501646 538634
rect 501882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 64826 534454
rect 65062 534218 65146 534454
rect 65382 534218 100826 534454
rect 101062 534218 101146 534454
rect 101382 534218 136826 534454
rect 137062 534218 137146 534454
rect 137382 534218 172826 534454
rect 173062 534218 173146 534454
rect 173382 534218 208826 534454
rect 209062 534218 209146 534454
rect 209382 534218 244826 534454
rect 245062 534218 245146 534454
rect 245382 534218 280826 534454
rect 281062 534218 281146 534454
rect 281382 534218 316826 534454
rect 317062 534218 317146 534454
rect 317382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 388826 534454
rect 389062 534218 389146 534454
rect 389382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 496826 534454
rect 497062 534218 497146 534454
rect 497382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 64826 534134
rect 65062 533898 65146 534134
rect 65382 533898 100826 534134
rect 101062 533898 101146 534134
rect 101382 533898 136826 534134
rect 137062 533898 137146 534134
rect 137382 533898 172826 534134
rect 173062 533898 173146 534134
rect 173382 533898 208826 534134
rect 209062 533898 209146 534134
rect 209382 533898 244826 534134
rect 245062 533898 245146 534134
rect 245382 533898 280826 534134
rect 281062 533898 281146 534134
rect 281382 533898 316826 534134
rect 317062 533898 317146 534134
rect 317382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 388826 534134
rect 389062 533898 389146 534134
rect 389382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 496826 534134
rect 497062 533898 497146 534134
rect 497382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 60326 529954
rect 60562 529718 60646 529954
rect 60882 529718 96326 529954
rect 96562 529718 96646 529954
rect 96882 529718 132326 529954
rect 132562 529718 132646 529954
rect 132882 529718 168326 529954
rect 168562 529718 168646 529954
rect 168882 529718 204326 529954
rect 204562 529718 204646 529954
rect 204882 529718 240326 529954
rect 240562 529718 240646 529954
rect 240882 529718 276326 529954
rect 276562 529718 276646 529954
rect 276882 529718 312326 529954
rect 312562 529718 312646 529954
rect 312882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 384326 529954
rect 384562 529718 384646 529954
rect 384882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 492326 529954
rect 492562 529718 492646 529954
rect 492882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 60326 529634
rect 60562 529398 60646 529634
rect 60882 529398 96326 529634
rect 96562 529398 96646 529634
rect 96882 529398 132326 529634
rect 132562 529398 132646 529634
rect 132882 529398 168326 529634
rect 168562 529398 168646 529634
rect 168882 529398 204326 529634
rect 204562 529398 204646 529634
rect 204882 529398 240326 529634
rect 240562 529398 240646 529634
rect 240882 529398 276326 529634
rect 276562 529398 276646 529634
rect 276882 529398 312326 529634
rect 312562 529398 312646 529634
rect 312882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 384326 529634
rect 384562 529398 384646 529634
rect 384882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 492326 529634
rect 492562 529398 492646 529634
rect 492882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 51326 520954
rect 51562 520718 51646 520954
rect 51882 520718 87326 520954
rect 87562 520718 87646 520954
rect 87882 520718 123326 520954
rect 123562 520718 123646 520954
rect 123882 520718 159326 520954
rect 159562 520718 159646 520954
rect 159882 520718 195326 520954
rect 195562 520718 195646 520954
rect 195882 520718 231326 520954
rect 231562 520718 231646 520954
rect 231882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 303326 520954
rect 303562 520718 303646 520954
rect 303882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 375326 520954
rect 375562 520718 375646 520954
rect 375882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 483326 520954
rect 483562 520718 483646 520954
rect 483882 520718 519326 520954
rect 519562 520718 519646 520954
rect 519882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 51326 520634
rect 51562 520398 51646 520634
rect 51882 520398 87326 520634
rect 87562 520398 87646 520634
rect 87882 520398 123326 520634
rect 123562 520398 123646 520634
rect 123882 520398 159326 520634
rect 159562 520398 159646 520634
rect 159882 520398 195326 520634
rect 195562 520398 195646 520634
rect 195882 520398 231326 520634
rect 231562 520398 231646 520634
rect 231882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 303326 520634
rect 303562 520398 303646 520634
rect 303882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 375326 520634
rect 375562 520398 375646 520634
rect 375882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 483326 520634
rect 483562 520398 483646 520634
rect 483882 520398 519326 520634
rect 519562 520398 519646 520634
rect 519882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 82826 516454
rect 83062 516218 83146 516454
rect 83382 516218 118826 516454
rect 119062 516218 119146 516454
rect 119382 516218 154826 516454
rect 155062 516218 155146 516454
rect 155382 516218 190826 516454
rect 191062 516218 191146 516454
rect 191382 516218 226826 516454
rect 227062 516218 227146 516454
rect 227382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 298826 516454
rect 299062 516218 299146 516454
rect 299382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 370826 516454
rect 371062 516218 371146 516454
rect 371382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 478826 516454
rect 479062 516218 479146 516454
rect 479382 516218 514826 516454
rect 515062 516218 515146 516454
rect 515382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 82826 516134
rect 83062 515898 83146 516134
rect 83382 515898 118826 516134
rect 119062 515898 119146 516134
rect 119382 515898 154826 516134
rect 155062 515898 155146 516134
rect 155382 515898 190826 516134
rect 191062 515898 191146 516134
rect 191382 515898 226826 516134
rect 227062 515898 227146 516134
rect 227382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 298826 516134
rect 299062 515898 299146 516134
rect 299382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 370826 516134
rect 371062 515898 371146 516134
rect 371382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 478826 516134
rect 479062 515898 479146 516134
rect 479382 515898 514826 516134
rect 515062 515898 515146 516134
rect 515382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 78326 511954
rect 78562 511718 78646 511954
rect 78882 511718 114326 511954
rect 114562 511718 114646 511954
rect 114882 511718 150326 511954
rect 150562 511718 150646 511954
rect 150882 511718 186326 511954
rect 186562 511718 186646 511954
rect 186882 511718 222326 511954
rect 222562 511718 222646 511954
rect 222882 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 294326 511954
rect 294562 511718 294646 511954
rect 294882 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 366326 511954
rect 366562 511718 366646 511954
rect 366882 511718 402326 511954
rect 402562 511718 402646 511954
rect 402882 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 510326 511954
rect 510562 511718 510646 511954
rect 510882 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 78326 511634
rect 78562 511398 78646 511634
rect 78882 511398 114326 511634
rect 114562 511398 114646 511634
rect 114882 511398 150326 511634
rect 150562 511398 150646 511634
rect 150882 511398 186326 511634
rect 186562 511398 186646 511634
rect 186882 511398 222326 511634
rect 222562 511398 222646 511634
rect 222882 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 294326 511634
rect 294562 511398 294646 511634
rect 294882 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 366326 511634
rect 366562 511398 366646 511634
rect 366882 511398 402326 511634
rect 402562 511398 402646 511634
rect 402882 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 510326 511634
rect 510562 511398 510646 511634
rect 510882 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 69326 502954
rect 69562 502718 69646 502954
rect 69882 502718 105326 502954
rect 105562 502718 105646 502954
rect 105882 502718 141326 502954
rect 141562 502718 141646 502954
rect 141882 502718 177326 502954
rect 177562 502718 177646 502954
rect 177882 502718 213326 502954
rect 213562 502718 213646 502954
rect 213882 502718 249326 502954
rect 249562 502718 249646 502954
rect 249882 502718 285326 502954
rect 285562 502718 285646 502954
rect 285882 502718 321326 502954
rect 321562 502718 321646 502954
rect 321882 502718 357326 502954
rect 357562 502718 357646 502954
rect 357882 502718 393326 502954
rect 393562 502718 393646 502954
rect 393882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 501326 502954
rect 501562 502718 501646 502954
rect 501882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 69326 502634
rect 69562 502398 69646 502634
rect 69882 502398 105326 502634
rect 105562 502398 105646 502634
rect 105882 502398 141326 502634
rect 141562 502398 141646 502634
rect 141882 502398 177326 502634
rect 177562 502398 177646 502634
rect 177882 502398 213326 502634
rect 213562 502398 213646 502634
rect 213882 502398 249326 502634
rect 249562 502398 249646 502634
rect 249882 502398 285326 502634
rect 285562 502398 285646 502634
rect 285882 502398 321326 502634
rect 321562 502398 321646 502634
rect 321882 502398 357326 502634
rect 357562 502398 357646 502634
rect 357882 502398 393326 502634
rect 393562 502398 393646 502634
rect 393882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 501326 502634
rect 501562 502398 501646 502634
rect 501882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 64826 498454
rect 65062 498218 65146 498454
rect 65382 498218 100826 498454
rect 101062 498218 101146 498454
rect 101382 498218 136826 498454
rect 137062 498218 137146 498454
rect 137382 498218 172826 498454
rect 173062 498218 173146 498454
rect 173382 498218 208826 498454
rect 209062 498218 209146 498454
rect 209382 498218 244826 498454
rect 245062 498218 245146 498454
rect 245382 498218 280826 498454
rect 281062 498218 281146 498454
rect 281382 498218 316826 498454
rect 317062 498218 317146 498454
rect 317382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 388826 498454
rect 389062 498218 389146 498454
rect 389382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 496826 498454
rect 497062 498218 497146 498454
rect 497382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 64826 498134
rect 65062 497898 65146 498134
rect 65382 497898 100826 498134
rect 101062 497898 101146 498134
rect 101382 497898 136826 498134
rect 137062 497898 137146 498134
rect 137382 497898 172826 498134
rect 173062 497898 173146 498134
rect 173382 497898 208826 498134
rect 209062 497898 209146 498134
rect 209382 497898 244826 498134
rect 245062 497898 245146 498134
rect 245382 497898 280826 498134
rect 281062 497898 281146 498134
rect 281382 497898 316826 498134
rect 317062 497898 317146 498134
rect 317382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 388826 498134
rect 389062 497898 389146 498134
rect 389382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 496826 498134
rect 497062 497898 497146 498134
rect 497382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 60326 493954
rect 60562 493718 60646 493954
rect 60882 493718 96326 493954
rect 96562 493718 96646 493954
rect 96882 493718 132326 493954
rect 132562 493718 132646 493954
rect 132882 493718 168326 493954
rect 168562 493718 168646 493954
rect 168882 493718 204326 493954
rect 204562 493718 204646 493954
rect 204882 493718 240326 493954
rect 240562 493718 240646 493954
rect 240882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 60326 493634
rect 60562 493398 60646 493634
rect 60882 493398 96326 493634
rect 96562 493398 96646 493634
rect 96882 493398 132326 493634
rect 132562 493398 132646 493634
rect 132882 493398 168326 493634
rect 168562 493398 168646 493634
rect 168882 493398 204326 493634
rect 204562 493398 204646 493634
rect 204882 493398 240326 493634
rect 240562 493398 240646 493634
rect 240882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 51326 484954
rect 51562 484718 51646 484954
rect 51882 484718 87326 484954
rect 87562 484718 87646 484954
rect 87882 484718 123326 484954
rect 123562 484718 123646 484954
rect 123882 484718 159326 484954
rect 159562 484718 159646 484954
rect 159882 484718 195326 484954
rect 195562 484718 195646 484954
rect 195882 484718 231326 484954
rect 231562 484718 231646 484954
rect 231882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 51326 484634
rect 51562 484398 51646 484634
rect 51882 484398 87326 484634
rect 87562 484398 87646 484634
rect 87882 484398 123326 484634
rect 123562 484398 123646 484634
rect 123882 484398 159326 484634
rect 159562 484398 159646 484634
rect 159882 484398 195326 484634
rect 195562 484398 195646 484634
rect 195882 484398 231326 484634
rect 231562 484398 231646 484634
rect 231882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 82826 480454
rect 83062 480218 83146 480454
rect 83382 480218 118826 480454
rect 119062 480218 119146 480454
rect 119382 480218 154826 480454
rect 155062 480218 155146 480454
rect 155382 480218 190826 480454
rect 191062 480218 191146 480454
rect 191382 480218 226826 480454
rect 227062 480218 227146 480454
rect 227382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 82826 480134
rect 83062 479898 83146 480134
rect 83382 479898 118826 480134
rect 119062 479898 119146 480134
rect 119382 479898 154826 480134
rect 155062 479898 155146 480134
rect 155382 479898 190826 480134
rect 191062 479898 191146 480134
rect 191382 479898 226826 480134
rect 227062 479898 227146 480134
rect 227382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 78326 475954
rect 78562 475718 78646 475954
rect 78882 475718 114326 475954
rect 114562 475718 114646 475954
rect 114882 475718 150326 475954
rect 150562 475718 150646 475954
rect 150882 475718 186326 475954
rect 186562 475718 186646 475954
rect 186882 475718 222326 475954
rect 222562 475718 222646 475954
rect 222882 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 78326 475634
rect 78562 475398 78646 475634
rect 78882 475398 114326 475634
rect 114562 475398 114646 475634
rect 114882 475398 150326 475634
rect 150562 475398 150646 475634
rect 150882 475398 186326 475634
rect 186562 475398 186646 475634
rect 186882 475398 222326 475634
rect 222562 475398 222646 475634
rect 222882 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 69326 466954
rect 69562 466718 69646 466954
rect 69882 466718 105326 466954
rect 105562 466718 105646 466954
rect 105882 466718 141326 466954
rect 141562 466718 141646 466954
rect 141882 466718 177326 466954
rect 177562 466718 177646 466954
rect 177882 466718 213326 466954
rect 213562 466718 213646 466954
rect 213882 466718 249326 466954
rect 249562 466718 249646 466954
rect 249882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 69326 466634
rect 69562 466398 69646 466634
rect 69882 466398 105326 466634
rect 105562 466398 105646 466634
rect 105882 466398 141326 466634
rect 141562 466398 141646 466634
rect 141882 466398 177326 466634
rect 177562 466398 177646 466634
rect 177882 466398 213326 466634
rect 213562 466398 213646 466634
rect 213882 466398 249326 466634
rect 249562 466398 249646 466634
rect 249882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 64826 462454
rect 65062 462218 65146 462454
rect 65382 462218 100826 462454
rect 101062 462218 101146 462454
rect 101382 462218 136826 462454
rect 137062 462218 137146 462454
rect 137382 462218 172826 462454
rect 173062 462218 173146 462454
rect 173382 462218 208826 462454
rect 209062 462218 209146 462454
rect 209382 462218 244826 462454
rect 245062 462218 245146 462454
rect 245382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 64826 462134
rect 65062 461898 65146 462134
rect 65382 461898 100826 462134
rect 101062 461898 101146 462134
rect 101382 461898 136826 462134
rect 137062 461898 137146 462134
rect 137382 461898 172826 462134
rect 173062 461898 173146 462134
rect 173382 461898 208826 462134
rect 209062 461898 209146 462134
rect 209382 461898 244826 462134
rect 245062 461898 245146 462134
rect 245382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 60326 457954
rect 60562 457718 60646 457954
rect 60882 457718 96326 457954
rect 96562 457718 96646 457954
rect 96882 457718 132326 457954
rect 132562 457718 132646 457954
rect 132882 457718 168326 457954
rect 168562 457718 168646 457954
rect 168882 457718 204326 457954
rect 204562 457718 204646 457954
rect 204882 457718 240326 457954
rect 240562 457718 240646 457954
rect 240882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 60326 457634
rect 60562 457398 60646 457634
rect 60882 457398 96326 457634
rect 96562 457398 96646 457634
rect 96882 457398 132326 457634
rect 132562 457398 132646 457634
rect 132882 457398 168326 457634
rect 168562 457398 168646 457634
rect 168882 457398 204326 457634
rect 204562 457398 204646 457634
rect 204882 457398 240326 457634
rect 240562 457398 240646 457634
rect 240882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 51326 448954
rect 51562 448718 51646 448954
rect 51882 448718 87326 448954
rect 87562 448718 87646 448954
rect 87882 448718 123326 448954
rect 123562 448718 123646 448954
rect 123882 448718 159326 448954
rect 159562 448718 159646 448954
rect 159882 448718 195326 448954
rect 195562 448718 195646 448954
rect 195882 448718 231326 448954
rect 231562 448718 231646 448954
rect 231882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 51326 448634
rect 51562 448398 51646 448634
rect 51882 448398 87326 448634
rect 87562 448398 87646 448634
rect 87882 448398 123326 448634
rect 123562 448398 123646 448634
rect 123882 448398 159326 448634
rect 159562 448398 159646 448634
rect 159882 448398 195326 448634
rect 195562 448398 195646 448634
rect 195882 448398 231326 448634
rect 231562 448398 231646 448634
rect 231882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 82826 444454
rect 83062 444218 83146 444454
rect 83382 444218 118826 444454
rect 119062 444218 119146 444454
rect 119382 444218 154826 444454
rect 155062 444218 155146 444454
rect 155382 444218 190826 444454
rect 191062 444218 191146 444454
rect 191382 444218 226826 444454
rect 227062 444218 227146 444454
rect 227382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 82826 444134
rect 83062 443898 83146 444134
rect 83382 443898 118826 444134
rect 119062 443898 119146 444134
rect 119382 443898 154826 444134
rect 155062 443898 155146 444134
rect 155382 443898 190826 444134
rect 191062 443898 191146 444134
rect 191382 443898 226826 444134
rect 227062 443898 227146 444134
rect 227382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 78326 439954
rect 78562 439718 78646 439954
rect 78882 439718 114326 439954
rect 114562 439718 114646 439954
rect 114882 439718 150326 439954
rect 150562 439718 150646 439954
rect 150882 439718 186326 439954
rect 186562 439718 186646 439954
rect 186882 439718 222326 439954
rect 222562 439718 222646 439954
rect 222882 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 78326 439634
rect 78562 439398 78646 439634
rect 78882 439398 114326 439634
rect 114562 439398 114646 439634
rect 114882 439398 150326 439634
rect 150562 439398 150646 439634
rect 150882 439398 186326 439634
rect 186562 439398 186646 439634
rect 186882 439398 222326 439634
rect 222562 439398 222646 439634
rect 222882 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 69326 430954
rect 69562 430718 69646 430954
rect 69882 430718 105326 430954
rect 105562 430718 105646 430954
rect 105882 430718 141326 430954
rect 141562 430718 141646 430954
rect 141882 430718 177326 430954
rect 177562 430718 177646 430954
rect 177882 430718 213326 430954
rect 213562 430718 213646 430954
rect 213882 430718 249326 430954
rect 249562 430718 249646 430954
rect 249882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 69326 430634
rect 69562 430398 69646 430634
rect 69882 430398 105326 430634
rect 105562 430398 105646 430634
rect 105882 430398 141326 430634
rect 141562 430398 141646 430634
rect 141882 430398 177326 430634
rect 177562 430398 177646 430634
rect 177882 430398 213326 430634
rect 213562 430398 213646 430634
rect 213882 430398 249326 430634
rect 249562 430398 249646 430634
rect 249882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 64826 426454
rect 65062 426218 65146 426454
rect 65382 426218 100826 426454
rect 101062 426218 101146 426454
rect 101382 426218 136826 426454
rect 137062 426218 137146 426454
rect 137382 426218 172826 426454
rect 173062 426218 173146 426454
rect 173382 426218 208826 426454
rect 209062 426218 209146 426454
rect 209382 426218 244826 426454
rect 245062 426218 245146 426454
rect 245382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 64826 426134
rect 65062 425898 65146 426134
rect 65382 425898 100826 426134
rect 101062 425898 101146 426134
rect 101382 425898 136826 426134
rect 137062 425898 137146 426134
rect 137382 425898 172826 426134
rect 173062 425898 173146 426134
rect 173382 425898 208826 426134
rect 209062 425898 209146 426134
rect 209382 425898 244826 426134
rect 245062 425898 245146 426134
rect 245382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 60326 421954
rect 60562 421718 60646 421954
rect 60882 421718 96326 421954
rect 96562 421718 96646 421954
rect 96882 421718 132326 421954
rect 132562 421718 132646 421954
rect 132882 421718 168326 421954
rect 168562 421718 168646 421954
rect 168882 421718 204326 421954
rect 204562 421718 204646 421954
rect 204882 421718 240326 421954
rect 240562 421718 240646 421954
rect 240882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 60326 421634
rect 60562 421398 60646 421634
rect 60882 421398 96326 421634
rect 96562 421398 96646 421634
rect 96882 421398 132326 421634
rect 132562 421398 132646 421634
rect 132882 421398 168326 421634
rect 168562 421398 168646 421634
rect 168882 421398 204326 421634
rect 204562 421398 204646 421634
rect 204882 421398 240326 421634
rect 240562 421398 240646 421634
rect 240882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 51326 412954
rect 51562 412718 51646 412954
rect 51882 412718 87326 412954
rect 87562 412718 87646 412954
rect 87882 412718 123326 412954
rect 123562 412718 123646 412954
rect 123882 412718 159326 412954
rect 159562 412718 159646 412954
rect 159882 412718 195326 412954
rect 195562 412718 195646 412954
rect 195882 412718 231326 412954
rect 231562 412718 231646 412954
rect 231882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 51326 412634
rect 51562 412398 51646 412634
rect 51882 412398 87326 412634
rect 87562 412398 87646 412634
rect 87882 412398 123326 412634
rect 123562 412398 123646 412634
rect 123882 412398 159326 412634
rect 159562 412398 159646 412634
rect 159882 412398 195326 412634
rect 195562 412398 195646 412634
rect 195882 412398 231326 412634
rect 231562 412398 231646 412634
rect 231882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 82826 408454
rect 83062 408218 83146 408454
rect 83382 408218 118826 408454
rect 119062 408218 119146 408454
rect 119382 408218 154826 408454
rect 155062 408218 155146 408454
rect 155382 408218 190826 408454
rect 191062 408218 191146 408454
rect 191382 408218 226826 408454
rect 227062 408218 227146 408454
rect 227382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 82826 408134
rect 83062 407898 83146 408134
rect 83382 407898 118826 408134
rect 119062 407898 119146 408134
rect 119382 407898 154826 408134
rect 155062 407898 155146 408134
rect 155382 407898 190826 408134
rect 191062 407898 191146 408134
rect 191382 407898 226826 408134
rect 227062 407898 227146 408134
rect 227382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 78326 403954
rect 78562 403718 78646 403954
rect 78882 403718 114326 403954
rect 114562 403718 114646 403954
rect 114882 403718 150326 403954
rect 150562 403718 150646 403954
rect 150882 403718 186326 403954
rect 186562 403718 186646 403954
rect 186882 403718 222326 403954
rect 222562 403718 222646 403954
rect 222882 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 78326 403634
rect 78562 403398 78646 403634
rect 78882 403398 114326 403634
rect 114562 403398 114646 403634
rect 114882 403398 150326 403634
rect 150562 403398 150646 403634
rect 150882 403398 186326 403634
rect 186562 403398 186646 403634
rect 186882 403398 222326 403634
rect 222562 403398 222646 403634
rect 222882 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 69326 394954
rect 69562 394718 69646 394954
rect 69882 394718 105326 394954
rect 105562 394718 105646 394954
rect 105882 394718 141326 394954
rect 141562 394718 141646 394954
rect 141882 394718 177326 394954
rect 177562 394718 177646 394954
rect 177882 394718 213326 394954
rect 213562 394718 213646 394954
rect 213882 394718 249326 394954
rect 249562 394718 249646 394954
rect 249882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 69326 394634
rect 69562 394398 69646 394634
rect 69882 394398 105326 394634
rect 105562 394398 105646 394634
rect 105882 394398 141326 394634
rect 141562 394398 141646 394634
rect 141882 394398 177326 394634
rect 177562 394398 177646 394634
rect 177882 394398 213326 394634
rect 213562 394398 213646 394634
rect 213882 394398 249326 394634
rect 249562 394398 249646 394634
rect 249882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 64826 390454
rect 65062 390218 65146 390454
rect 65382 390218 100826 390454
rect 101062 390218 101146 390454
rect 101382 390218 136826 390454
rect 137062 390218 137146 390454
rect 137382 390218 172826 390454
rect 173062 390218 173146 390454
rect 173382 390218 208826 390454
rect 209062 390218 209146 390454
rect 209382 390218 244826 390454
rect 245062 390218 245146 390454
rect 245382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 64826 390134
rect 65062 389898 65146 390134
rect 65382 389898 100826 390134
rect 101062 389898 101146 390134
rect 101382 389898 136826 390134
rect 137062 389898 137146 390134
rect 137382 389898 172826 390134
rect 173062 389898 173146 390134
rect 173382 389898 208826 390134
rect 209062 389898 209146 390134
rect 209382 389898 244826 390134
rect 245062 389898 245146 390134
rect 245382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 60326 385954
rect 60562 385718 60646 385954
rect 60882 385718 96326 385954
rect 96562 385718 96646 385954
rect 96882 385718 132326 385954
rect 132562 385718 132646 385954
rect 132882 385718 168326 385954
rect 168562 385718 168646 385954
rect 168882 385718 204326 385954
rect 204562 385718 204646 385954
rect 204882 385718 240326 385954
rect 240562 385718 240646 385954
rect 240882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 60326 385634
rect 60562 385398 60646 385634
rect 60882 385398 96326 385634
rect 96562 385398 96646 385634
rect 96882 385398 132326 385634
rect 132562 385398 132646 385634
rect 132882 385398 168326 385634
rect 168562 385398 168646 385634
rect 168882 385398 204326 385634
rect 204562 385398 204646 385634
rect 204882 385398 240326 385634
rect 240562 385398 240646 385634
rect 240882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 51326 376954
rect 51562 376718 51646 376954
rect 51882 376718 87326 376954
rect 87562 376718 87646 376954
rect 87882 376718 123326 376954
rect 123562 376718 123646 376954
rect 123882 376718 159326 376954
rect 159562 376718 159646 376954
rect 159882 376718 195326 376954
rect 195562 376718 195646 376954
rect 195882 376718 231326 376954
rect 231562 376718 231646 376954
rect 231882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 51326 376634
rect 51562 376398 51646 376634
rect 51882 376398 87326 376634
rect 87562 376398 87646 376634
rect 87882 376398 123326 376634
rect 123562 376398 123646 376634
rect 123882 376398 159326 376634
rect 159562 376398 159646 376634
rect 159882 376398 195326 376634
rect 195562 376398 195646 376634
rect 195882 376398 231326 376634
rect 231562 376398 231646 376634
rect 231882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 82826 372454
rect 83062 372218 83146 372454
rect 83382 372218 118826 372454
rect 119062 372218 119146 372454
rect 119382 372218 154826 372454
rect 155062 372218 155146 372454
rect 155382 372218 190826 372454
rect 191062 372218 191146 372454
rect 191382 372218 226826 372454
rect 227062 372218 227146 372454
rect 227382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 82826 372134
rect 83062 371898 83146 372134
rect 83382 371898 118826 372134
rect 119062 371898 119146 372134
rect 119382 371898 154826 372134
rect 155062 371898 155146 372134
rect 155382 371898 190826 372134
rect 191062 371898 191146 372134
rect 191382 371898 226826 372134
rect 227062 371898 227146 372134
rect 227382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 78326 367954
rect 78562 367718 78646 367954
rect 78882 367718 114326 367954
rect 114562 367718 114646 367954
rect 114882 367718 150326 367954
rect 150562 367718 150646 367954
rect 150882 367718 186326 367954
rect 186562 367718 186646 367954
rect 186882 367718 222326 367954
rect 222562 367718 222646 367954
rect 222882 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 78326 367634
rect 78562 367398 78646 367634
rect 78882 367398 114326 367634
rect 114562 367398 114646 367634
rect 114882 367398 150326 367634
rect 150562 367398 150646 367634
rect 150882 367398 186326 367634
rect 186562 367398 186646 367634
rect 186882 367398 222326 367634
rect 222562 367398 222646 367634
rect 222882 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 69326 358954
rect 69562 358718 69646 358954
rect 69882 358718 105326 358954
rect 105562 358718 105646 358954
rect 105882 358718 141326 358954
rect 141562 358718 141646 358954
rect 141882 358718 177326 358954
rect 177562 358718 177646 358954
rect 177882 358718 213326 358954
rect 213562 358718 213646 358954
rect 213882 358718 249326 358954
rect 249562 358718 249646 358954
rect 249882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 69326 358634
rect 69562 358398 69646 358634
rect 69882 358398 105326 358634
rect 105562 358398 105646 358634
rect 105882 358398 141326 358634
rect 141562 358398 141646 358634
rect 141882 358398 177326 358634
rect 177562 358398 177646 358634
rect 177882 358398 213326 358634
rect 213562 358398 213646 358634
rect 213882 358398 249326 358634
rect 249562 358398 249646 358634
rect 249882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 64826 354454
rect 65062 354218 65146 354454
rect 65382 354218 100826 354454
rect 101062 354218 101146 354454
rect 101382 354218 136826 354454
rect 137062 354218 137146 354454
rect 137382 354218 172826 354454
rect 173062 354218 173146 354454
rect 173382 354218 208826 354454
rect 209062 354218 209146 354454
rect 209382 354218 244826 354454
rect 245062 354218 245146 354454
rect 245382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 64826 354134
rect 65062 353898 65146 354134
rect 65382 353898 100826 354134
rect 101062 353898 101146 354134
rect 101382 353898 136826 354134
rect 137062 353898 137146 354134
rect 137382 353898 172826 354134
rect 173062 353898 173146 354134
rect 173382 353898 208826 354134
rect 209062 353898 209146 354134
rect 209382 353898 244826 354134
rect 245062 353898 245146 354134
rect 245382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 60326 349954
rect 60562 349718 60646 349954
rect 60882 349718 96326 349954
rect 96562 349718 96646 349954
rect 96882 349718 132326 349954
rect 132562 349718 132646 349954
rect 132882 349718 168326 349954
rect 168562 349718 168646 349954
rect 168882 349718 204326 349954
rect 204562 349718 204646 349954
rect 204882 349718 240326 349954
rect 240562 349718 240646 349954
rect 240882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 60326 349634
rect 60562 349398 60646 349634
rect 60882 349398 96326 349634
rect 96562 349398 96646 349634
rect 96882 349398 132326 349634
rect 132562 349398 132646 349634
rect 132882 349398 168326 349634
rect 168562 349398 168646 349634
rect 168882 349398 204326 349634
rect 204562 349398 204646 349634
rect 204882 349398 240326 349634
rect 240562 349398 240646 349634
rect 240882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 51326 340954
rect 51562 340718 51646 340954
rect 51882 340718 87326 340954
rect 87562 340718 87646 340954
rect 87882 340718 123326 340954
rect 123562 340718 123646 340954
rect 123882 340718 159326 340954
rect 159562 340718 159646 340954
rect 159882 340718 195326 340954
rect 195562 340718 195646 340954
rect 195882 340718 231326 340954
rect 231562 340718 231646 340954
rect 231882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 51326 340634
rect 51562 340398 51646 340634
rect 51882 340398 87326 340634
rect 87562 340398 87646 340634
rect 87882 340398 123326 340634
rect 123562 340398 123646 340634
rect 123882 340398 159326 340634
rect 159562 340398 159646 340634
rect 159882 340398 195326 340634
rect 195562 340398 195646 340634
rect 195882 340398 231326 340634
rect 231562 340398 231646 340634
rect 231882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 82826 336454
rect 83062 336218 83146 336454
rect 83382 336218 118826 336454
rect 119062 336218 119146 336454
rect 119382 336218 154826 336454
rect 155062 336218 155146 336454
rect 155382 336218 190826 336454
rect 191062 336218 191146 336454
rect 191382 336218 226826 336454
rect 227062 336218 227146 336454
rect 227382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 82826 336134
rect 83062 335898 83146 336134
rect 83382 335898 118826 336134
rect 119062 335898 119146 336134
rect 119382 335898 154826 336134
rect 155062 335898 155146 336134
rect 155382 335898 190826 336134
rect 191062 335898 191146 336134
rect 191382 335898 226826 336134
rect 227062 335898 227146 336134
rect 227382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 78326 331954
rect 78562 331718 78646 331954
rect 78882 331718 114326 331954
rect 114562 331718 114646 331954
rect 114882 331718 150326 331954
rect 150562 331718 150646 331954
rect 150882 331718 186326 331954
rect 186562 331718 186646 331954
rect 186882 331718 222326 331954
rect 222562 331718 222646 331954
rect 222882 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 330326 331954
rect 330562 331718 330646 331954
rect 330882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 78326 331634
rect 78562 331398 78646 331634
rect 78882 331398 114326 331634
rect 114562 331398 114646 331634
rect 114882 331398 150326 331634
rect 150562 331398 150646 331634
rect 150882 331398 186326 331634
rect 186562 331398 186646 331634
rect 186882 331398 222326 331634
rect 222562 331398 222646 331634
rect 222882 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 330326 331634
rect 330562 331398 330646 331634
rect 330882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 69326 322954
rect 69562 322718 69646 322954
rect 69882 322718 105326 322954
rect 105562 322718 105646 322954
rect 105882 322718 141326 322954
rect 141562 322718 141646 322954
rect 141882 322718 177326 322954
rect 177562 322718 177646 322954
rect 177882 322718 213326 322954
rect 213562 322718 213646 322954
rect 213882 322718 249326 322954
rect 249562 322718 249646 322954
rect 249882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 321326 322954
rect 321562 322718 321646 322954
rect 321882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 69326 322634
rect 69562 322398 69646 322634
rect 69882 322398 105326 322634
rect 105562 322398 105646 322634
rect 105882 322398 141326 322634
rect 141562 322398 141646 322634
rect 141882 322398 177326 322634
rect 177562 322398 177646 322634
rect 177882 322398 213326 322634
rect 213562 322398 213646 322634
rect 213882 322398 249326 322634
rect 249562 322398 249646 322634
rect 249882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 321326 322634
rect 321562 322398 321646 322634
rect 321882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 64826 318454
rect 65062 318218 65146 318454
rect 65382 318218 100826 318454
rect 101062 318218 101146 318454
rect 101382 318218 136826 318454
rect 137062 318218 137146 318454
rect 137382 318218 172826 318454
rect 173062 318218 173146 318454
rect 173382 318218 208826 318454
rect 209062 318218 209146 318454
rect 209382 318218 244826 318454
rect 245062 318218 245146 318454
rect 245382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 316826 318454
rect 317062 318218 317146 318454
rect 317382 318218 352826 318454
rect 353062 318218 353146 318454
rect 353382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 64826 318134
rect 65062 317898 65146 318134
rect 65382 317898 100826 318134
rect 101062 317898 101146 318134
rect 101382 317898 136826 318134
rect 137062 317898 137146 318134
rect 137382 317898 172826 318134
rect 173062 317898 173146 318134
rect 173382 317898 208826 318134
rect 209062 317898 209146 318134
rect 209382 317898 244826 318134
rect 245062 317898 245146 318134
rect 245382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 316826 318134
rect 317062 317898 317146 318134
rect 317382 317898 352826 318134
rect 353062 317898 353146 318134
rect 353382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 60326 313954
rect 60562 313718 60646 313954
rect 60882 313718 96326 313954
rect 96562 313718 96646 313954
rect 96882 313718 132326 313954
rect 132562 313718 132646 313954
rect 132882 313718 168326 313954
rect 168562 313718 168646 313954
rect 168882 313718 204326 313954
rect 204562 313718 204646 313954
rect 204882 313718 240326 313954
rect 240562 313718 240646 313954
rect 240882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 312326 313954
rect 312562 313718 312646 313954
rect 312882 313718 348326 313954
rect 348562 313718 348646 313954
rect 348882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 60326 313634
rect 60562 313398 60646 313634
rect 60882 313398 96326 313634
rect 96562 313398 96646 313634
rect 96882 313398 132326 313634
rect 132562 313398 132646 313634
rect 132882 313398 168326 313634
rect 168562 313398 168646 313634
rect 168882 313398 204326 313634
rect 204562 313398 204646 313634
rect 204882 313398 240326 313634
rect 240562 313398 240646 313634
rect 240882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 312326 313634
rect 312562 313398 312646 313634
rect 312882 313398 348326 313634
rect 348562 313398 348646 313634
rect 348882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 51326 304954
rect 51562 304718 51646 304954
rect 51882 304718 87326 304954
rect 87562 304718 87646 304954
rect 87882 304718 123326 304954
rect 123562 304718 123646 304954
rect 123882 304718 159326 304954
rect 159562 304718 159646 304954
rect 159882 304718 195326 304954
rect 195562 304718 195646 304954
rect 195882 304718 231326 304954
rect 231562 304718 231646 304954
rect 231882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 303326 304954
rect 303562 304718 303646 304954
rect 303882 304718 339326 304954
rect 339562 304718 339646 304954
rect 339882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 51326 304634
rect 51562 304398 51646 304634
rect 51882 304398 87326 304634
rect 87562 304398 87646 304634
rect 87882 304398 123326 304634
rect 123562 304398 123646 304634
rect 123882 304398 159326 304634
rect 159562 304398 159646 304634
rect 159882 304398 195326 304634
rect 195562 304398 195646 304634
rect 195882 304398 231326 304634
rect 231562 304398 231646 304634
rect 231882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 303326 304634
rect 303562 304398 303646 304634
rect 303882 304398 339326 304634
rect 339562 304398 339646 304634
rect 339882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 82826 300454
rect 83062 300218 83146 300454
rect 83382 300218 118826 300454
rect 119062 300218 119146 300454
rect 119382 300218 154826 300454
rect 155062 300218 155146 300454
rect 155382 300218 190826 300454
rect 191062 300218 191146 300454
rect 191382 300218 226826 300454
rect 227062 300218 227146 300454
rect 227382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 298826 300454
rect 299062 300218 299146 300454
rect 299382 300218 334826 300454
rect 335062 300218 335146 300454
rect 335382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 82826 300134
rect 83062 299898 83146 300134
rect 83382 299898 118826 300134
rect 119062 299898 119146 300134
rect 119382 299898 154826 300134
rect 155062 299898 155146 300134
rect 155382 299898 190826 300134
rect 191062 299898 191146 300134
rect 191382 299898 226826 300134
rect 227062 299898 227146 300134
rect 227382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 298826 300134
rect 299062 299898 299146 300134
rect 299382 299898 334826 300134
rect 335062 299898 335146 300134
rect 335382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 78326 295954
rect 78562 295718 78646 295954
rect 78882 295718 114326 295954
rect 114562 295718 114646 295954
rect 114882 295718 150326 295954
rect 150562 295718 150646 295954
rect 150882 295718 186326 295954
rect 186562 295718 186646 295954
rect 186882 295718 222326 295954
rect 222562 295718 222646 295954
rect 222882 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 330326 295954
rect 330562 295718 330646 295954
rect 330882 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 78326 295634
rect 78562 295398 78646 295634
rect 78882 295398 114326 295634
rect 114562 295398 114646 295634
rect 114882 295398 150326 295634
rect 150562 295398 150646 295634
rect 150882 295398 186326 295634
rect 186562 295398 186646 295634
rect 186882 295398 222326 295634
rect 222562 295398 222646 295634
rect 222882 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 330326 295634
rect 330562 295398 330646 295634
rect 330882 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 69326 286954
rect 69562 286718 69646 286954
rect 69882 286718 105326 286954
rect 105562 286718 105646 286954
rect 105882 286718 141326 286954
rect 141562 286718 141646 286954
rect 141882 286718 177326 286954
rect 177562 286718 177646 286954
rect 177882 286718 213326 286954
rect 213562 286718 213646 286954
rect 213882 286718 249326 286954
rect 249562 286718 249646 286954
rect 249882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 321326 286954
rect 321562 286718 321646 286954
rect 321882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 69326 286634
rect 69562 286398 69646 286634
rect 69882 286398 105326 286634
rect 105562 286398 105646 286634
rect 105882 286398 141326 286634
rect 141562 286398 141646 286634
rect 141882 286398 177326 286634
rect 177562 286398 177646 286634
rect 177882 286398 213326 286634
rect 213562 286398 213646 286634
rect 213882 286398 249326 286634
rect 249562 286398 249646 286634
rect 249882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 321326 286634
rect 321562 286398 321646 286634
rect 321882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 64826 282454
rect 65062 282218 65146 282454
rect 65382 282218 100826 282454
rect 101062 282218 101146 282454
rect 101382 282218 136826 282454
rect 137062 282218 137146 282454
rect 137382 282218 172826 282454
rect 173062 282218 173146 282454
rect 173382 282218 208826 282454
rect 209062 282218 209146 282454
rect 209382 282218 244826 282454
rect 245062 282218 245146 282454
rect 245382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 316826 282454
rect 317062 282218 317146 282454
rect 317382 282218 352826 282454
rect 353062 282218 353146 282454
rect 353382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 64826 282134
rect 65062 281898 65146 282134
rect 65382 281898 100826 282134
rect 101062 281898 101146 282134
rect 101382 281898 136826 282134
rect 137062 281898 137146 282134
rect 137382 281898 172826 282134
rect 173062 281898 173146 282134
rect 173382 281898 208826 282134
rect 209062 281898 209146 282134
rect 209382 281898 244826 282134
rect 245062 281898 245146 282134
rect 245382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 316826 282134
rect 317062 281898 317146 282134
rect 317382 281898 352826 282134
rect 353062 281898 353146 282134
rect 353382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 69326 250954
rect 69562 250718 69646 250954
rect 69882 250718 105326 250954
rect 105562 250718 105646 250954
rect 105882 250718 141326 250954
rect 141562 250718 141646 250954
rect 141882 250718 177326 250954
rect 177562 250718 177646 250954
rect 177882 250718 213326 250954
rect 213562 250718 213646 250954
rect 213882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 321326 250954
rect 321562 250718 321646 250954
rect 321882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 69326 250634
rect 69562 250398 69646 250634
rect 69882 250398 105326 250634
rect 105562 250398 105646 250634
rect 105882 250398 141326 250634
rect 141562 250398 141646 250634
rect 141882 250398 177326 250634
rect 177562 250398 177646 250634
rect 177882 250398 213326 250634
rect 213562 250398 213646 250634
rect 213882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 321326 250634
rect 321562 250398 321646 250634
rect 321882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 64826 246454
rect 65062 246218 65146 246454
rect 65382 246218 100826 246454
rect 101062 246218 101146 246454
rect 101382 246218 136826 246454
rect 137062 246218 137146 246454
rect 137382 246218 172826 246454
rect 173062 246218 173146 246454
rect 173382 246218 208826 246454
rect 209062 246218 209146 246454
rect 209382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 316826 246454
rect 317062 246218 317146 246454
rect 317382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 64826 246134
rect 65062 245898 65146 246134
rect 65382 245898 100826 246134
rect 101062 245898 101146 246134
rect 101382 245898 136826 246134
rect 137062 245898 137146 246134
rect 137382 245898 172826 246134
rect 173062 245898 173146 246134
rect 173382 245898 208826 246134
rect 209062 245898 209146 246134
rect 209382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 316826 246134
rect 317062 245898 317146 246134
rect 317382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 69326 214954
rect 69562 214718 69646 214954
rect 69882 214718 105326 214954
rect 105562 214718 105646 214954
rect 105882 214718 141326 214954
rect 141562 214718 141646 214954
rect 141882 214718 177326 214954
rect 177562 214718 177646 214954
rect 177882 214718 213326 214954
rect 213562 214718 213646 214954
rect 213882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 321326 214954
rect 321562 214718 321646 214954
rect 321882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 69326 214634
rect 69562 214398 69646 214634
rect 69882 214398 105326 214634
rect 105562 214398 105646 214634
rect 105882 214398 141326 214634
rect 141562 214398 141646 214634
rect 141882 214398 177326 214634
rect 177562 214398 177646 214634
rect 177882 214398 213326 214634
rect 213562 214398 213646 214634
rect 213882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 321326 214634
rect 321562 214398 321646 214634
rect 321882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 64826 210454
rect 65062 210218 65146 210454
rect 65382 210218 100826 210454
rect 101062 210218 101146 210454
rect 101382 210218 136826 210454
rect 137062 210218 137146 210454
rect 137382 210218 172826 210454
rect 173062 210218 173146 210454
rect 173382 210218 208826 210454
rect 209062 210218 209146 210454
rect 209382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 316826 210454
rect 317062 210218 317146 210454
rect 317382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 64826 210134
rect 65062 209898 65146 210134
rect 65382 209898 100826 210134
rect 101062 209898 101146 210134
rect 101382 209898 136826 210134
rect 137062 209898 137146 210134
rect 137382 209898 172826 210134
rect 173062 209898 173146 210134
rect 173382 209898 208826 210134
rect 209062 209898 209146 210134
rect 209382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 316826 210134
rect 317062 209898 317146 210134
rect 317382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 60326 205954
rect 60562 205718 60646 205954
rect 60882 205718 96326 205954
rect 96562 205718 96646 205954
rect 96882 205718 132326 205954
rect 132562 205718 132646 205954
rect 132882 205718 168326 205954
rect 168562 205718 168646 205954
rect 168882 205718 204326 205954
rect 204562 205718 204646 205954
rect 204882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 312326 205954
rect 312562 205718 312646 205954
rect 312882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 60326 205634
rect 60562 205398 60646 205634
rect 60882 205398 96326 205634
rect 96562 205398 96646 205634
rect 96882 205398 132326 205634
rect 132562 205398 132646 205634
rect 132882 205398 168326 205634
rect 168562 205398 168646 205634
rect 168882 205398 204326 205634
rect 204562 205398 204646 205634
rect 204882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 312326 205634
rect 312562 205398 312646 205634
rect 312882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 87326 196954
rect 87562 196718 87646 196954
rect 87882 196718 123326 196954
rect 123562 196718 123646 196954
rect 123882 196718 159326 196954
rect 159562 196718 159646 196954
rect 159882 196718 195326 196954
rect 195562 196718 195646 196954
rect 195882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 303326 196954
rect 303562 196718 303646 196954
rect 303882 196718 339326 196954
rect 339562 196718 339646 196954
rect 339882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 87326 196634
rect 87562 196398 87646 196634
rect 87882 196398 123326 196634
rect 123562 196398 123646 196634
rect 123882 196398 159326 196634
rect 159562 196398 159646 196634
rect 159882 196398 195326 196634
rect 195562 196398 195646 196634
rect 195882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 303326 196634
rect 303562 196398 303646 196634
rect 303882 196398 339326 196634
rect 339562 196398 339646 196634
rect 339882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 82826 192454
rect 83062 192218 83146 192454
rect 83382 192218 118826 192454
rect 119062 192218 119146 192454
rect 119382 192218 154826 192454
rect 155062 192218 155146 192454
rect 155382 192218 190826 192454
rect 191062 192218 191146 192454
rect 191382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 298826 192454
rect 299062 192218 299146 192454
rect 299382 192218 334826 192454
rect 335062 192218 335146 192454
rect 335382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 82826 192134
rect 83062 191898 83146 192134
rect 83382 191898 118826 192134
rect 119062 191898 119146 192134
rect 119382 191898 154826 192134
rect 155062 191898 155146 192134
rect 155382 191898 190826 192134
rect 191062 191898 191146 192134
rect 191382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 298826 192134
rect 299062 191898 299146 192134
rect 299382 191898 334826 192134
rect 335062 191898 335146 192134
rect 335382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 78326 187954
rect 78562 187718 78646 187954
rect 78882 187718 114326 187954
rect 114562 187718 114646 187954
rect 114882 187718 150326 187954
rect 150562 187718 150646 187954
rect 150882 187718 186326 187954
rect 186562 187718 186646 187954
rect 186882 187718 222326 187954
rect 222562 187718 222646 187954
rect 222882 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 330326 187954
rect 330562 187718 330646 187954
rect 330882 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 78326 187634
rect 78562 187398 78646 187634
rect 78882 187398 114326 187634
rect 114562 187398 114646 187634
rect 114882 187398 150326 187634
rect 150562 187398 150646 187634
rect 150882 187398 186326 187634
rect 186562 187398 186646 187634
rect 186882 187398 222326 187634
rect 222562 187398 222646 187634
rect 222882 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 330326 187634
rect 330562 187398 330646 187634
rect 330882 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 69326 178954
rect 69562 178718 69646 178954
rect 69882 178718 105326 178954
rect 105562 178718 105646 178954
rect 105882 178718 141326 178954
rect 141562 178718 141646 178954
rect 141882 178718 177326 178954
rect 177562 178718 177646 178954
rect 177882 178718 213326 178954
rect 213562 178718 213646 178954
rect 213882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 321326 178954
rect 321562 178718 321646 178954
rect 321882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 69326 178634
rect 69562 178398 69646 178634
rect 69882 178398 105326 178634
rect 105562 178398 105646 178634
rect 105882 178398 141326 178634
rect 141562 178398 141646 178634
rect 141882 178398 177326 178634
rect 177562 178398 177646 178634
rect 177882 178398 213326 178634
rect 213562 178398 213646 178634
rect 213882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 321326 178634
rect 321562 178398 321646 178634
rect 321882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 64826 174454
rect 65062 174218 65146 174454
rect 65382 174218 100826 174454
rect 101062 174218 101146 174454
rect 101382 174218 136826 174454
rect 137062 174218 137146 174454
rect 137382 174218 172826 174454
rect 173062 174218 173146 174454
rect 173382 174218 208826 174454
rect 209062 174218 209146 174454
rect 209382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 316826 174454
rect 317062 174218 317146 174454
rect 317382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 64826 174134
rect 65062 173898 65146 174134
rect 65382 173898 100826 174134
rect 101062 173898 101146 174134
rect 101382 173898 136826 174134
rect 137062 173898 137146 174134
rect 137382 173898 172826 174134
rect 173062 173898 173146 174134
rect 173382 173898 208826 174134
rect 209062 173898 209146 174134
rect 209382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 316826 174134
rect 317062 173898 317146 174134
rect 317382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 60326 169954
rect 60562 169718 60646 169954
rect 60882 169718 96326 169954
rect 96562 169718 96646 169954
rect 96882 169718 132326 169954
rect 132562 169718 132646 169954
rect 132882 169718 168326 169954
rect 168562 169718 168646 169954
rect 168882 169718 204326 169954
rect 204562 169718 204646 169954
rect 204882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 312326 169954
rect 312562 169718 312646 169954
rect 312882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 60326 169634
rect 60562 169398 60646 169634
rect 60882 169398 96326 169634
rect 96562 169398 96646 169634
rect 96882 169398 132326 169634
rect 132562 169398 132646 169634
rect 132882 169398 168326 169634
rect 168562 169398 168646 169634
rect 168882 169398 204326 169634
rect 204562 169398 204646 169634
rect 204882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 312326 169634
rect 312562 169398 312646 169634
rect 312882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 87326 160954
rect 87562 160718 87646 160954
rect 87882 160718 123326 160954
rect 123562 160718 123646 160954
rect 123882 160718 159326 160954
rect 159562 160718 159646 160954
rect 159882 160718 195326 160954
rect 195562 160718 195646 160954
rect 195882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 303326 160954
rect 303562 160718 303646 160954
rect 303882 160718 339326 160954
rect 339562 160718 339646 160954
rect 339882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 87326 160634
rect 87562 160398 87646 160634
rect 87882 160398 123326 160634
rect 123562 160398 123646 160634
rect 123882 160398 159326 160634
rect 159562 160398 159646 160634
rect 159882 160398 195326 160634
rect 195562 160398 195646 160634
rect 195882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 303326 160634
rect 303562 160398 303646 160634
rect 303882 160398 339326 160634
rect 339562 160398 339646 160634
rect 339882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 82826 156454
rect 83062 156218 83146 156454
rect 83382 156218 118826 156454
rect 119062 156218 119146 156454
rect 119382 156218 154826 156454
rect 155062 156218 155146 156454
rect 155382 156218 190826 156454
rect 191062 156218 191146 156454
rect 191382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 298826 156454
rect 299062 156218 299146 156454
rect 299382 156218 334826 156454
rect 335062 156218 335146 156454
rect 335382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 82826 156134
rect 83062 155898 83146 156134
rect 83382 155898 118826 156134
rect 119062 155898 119146 156134
rect 119382 155898 154826 156134
rect 155062 155898 155146 156134
rect 155382 155898 190826 156134
rect 191062 155898 191146 156134
rect 191382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 298826 156134
rect 299062 155898 299146 156134
rect 299382 155898 334826 156134
rect 335062 155898 335146 156134
rect 335382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 78326 151954
rect 78562 151718 78646 151954
rect 78882 151718 114326 151954
rect 114562 151718 114646 151954
rect 114882 151718 150326 151954
rect 150562 151718 150646 151954
rect 150882 151718 186326 151954
rect 186562 151718 186646 151954
rect 186882 151718 222326 151954
rect 222562 151718 222646 151954
rect 222882 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 330326 151954
rect 330562 151718 330646 151954
rect 330882 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 78326 151634
rect 78562 151398 78646 151634
rect 78882 151398 114326 151634
rect 114562 151398 114646 151634
rect 114882 151398 150326 151634
rect 150562 151398 150646 151634
rect 150882 151398 186326 151634
rect 186562 151398 186646 151634
rect 186882 151398 222326 151634
rect 222562 151398 222646 151634
rect 222882 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 330326 151634
rect 330562 151398 330646 151634
rect 330882 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 69326 142954
rect 69562 142718 69646 142954
rect 69882 142718 105326 142954
rect 105562 142718 105646 142954
rect 105882 142718 141326 142954
rect 141562 142718 141646 142954
rect 141882 142718 177326 142954
rect 177562 142718 177646 142954
rect 177882 142718 213326 142954
rect 213562 142718 213646 142954
rect 213882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 321326 142954
rect 321562 142718 321646 142954
rect 321882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 69326 142634
rect 69562 142398 69646 142634
rect 69882 142398 105326 142634
rect 105562 142398 105646 142634
rect 105882 142398 141326 142634
rect 141562 142398 141646 142634
rect 141882 142398 177326 142634
rect 177562 142398 177646 142634
rect 177882 142398 213326 142634
rect 213562 142398 213646 142634
rect 213882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 321326 142634
rect 321562 142398 321646 142634
rect 321882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 64826 138454
rect 65062 138218 65146 138454
rect 65382 138218 100826 138454
rect 101062 138218 101146 138454
rect 101382 138218 208826 138454
rect 209062 138218 209146 138454
rect 209382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 316826 138454
rect 317062 138218 317146 138454
rect 317382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 64826 138134
rect 65062 137898 65146 138134
rect 65382 137898 100826 138134
rect 101062 137898 101146 138134
rect 101382 137898 208826 138134
rect 209062 137898 209146 138134
rect 209382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 316826 138134
rect 317062 137898 317146 138134
rect 317382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 60326 133954
rect 60562 133718 60646 133954
rect 60882 133718 96326 133954
rect 96562 133718 96646 133954
rect 96882 133718 204326 133954
rect 204562 133718 204646 133954
rect 204882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 312326 133954
rect 312562 133718 312646 133954
rect 312882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 60326 133634
rect 60562 133398 60646 133634
rect 60882 133398 96326 133634
rect 96562 133398 96646 133634
rect 96882 133398 204326 133634
rect 204562 133398 204646 133634
rect 204882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 312326 133634
rect 312562 133398 312646 133634
rect 312882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 87326 124954
rect 87562 124718 87646 124954
rect 87882 124718 195326 124954
rect 195562 124718 195646 124954
rect 195882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 303326 124954
rect 303562 124718 303646 124954
rect 303882 124718 339326 124954
rect 339562 124718 339646 124954
rect 339882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 87326 124634
rect 87562 124398 87646 124634
rect 87882 124398 195326 124634
rect 195562 124398 195646 124634
rect 195882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 303326 124634
rect 303562 124398 303646 124634
rect 303882 124398 339326 124634
rect 339562 124398 339646 124634
rect 339882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 82826 120454
rect 83062 120218 83146 120454
rect 83382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 298826 120454
rect 299062 120218 299146 120454
rect 299382 120218 334826 120454
rect 335062 120218 335146 120454
rect 335382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 82826 120134
rect 83062 119898 83146 120134
rect 83382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 298826 120134
rect 299062 119898 299146 120134
rect 299382 119898 334826 120134
rect 335062 119898 335146 120134
rect 335382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 78326 115954
rect 78562 115718 78646 115954
rect 78882 115718 114326 115954
rect 114562 115718 114646 115954
rect 114882 115718 139610 115954
rect 139846 115718 170330 115954
rect 170566 115718 222326 115954
rect 222562 115718 222646 115954
rect 222882 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 330326 115954
rect 330562 115718 330646 115954
rect 330882 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 78326 115634
rect 78562 115398 78646 115634
rect 78882 115398 114326 115634
rect 114562 115398 114646 115634
rect 114882 115398 139610 115634
rect 139846 115398 170330 115634
rect 170566 115398 222326 115634
rect 222562 115398 222646 115634
rect 222882 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 330326 115634
rect 330562 115398 330646 115634
rect 330882 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 124250 111454
rect 124486 111218 154970 111454
rect 155206 111218 185690 111454
rect 185926 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 124250 111134
rect 124486 110898 154970 111134
rect 155206 110898 185690 111134
rect 185926 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 69326 106954
rect 69562 106718 69646 106954
rect 69882 106718 105326 106954
rect 105562 106718 105646 106954
rect 105882 106718 213326 106954
rect 213562 106718 213646 106954
rect 213882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 321326 106954
rect 321562 106718 321646 106954
rect 321882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 69326 106634
rect 69562 106398 69646 106634
rect 69882 106398 105326 106634
rect 105562 106398 105646 106634
rect 105882 106398 213326 106634
rect 213562 106398 213646 106634
rect 213882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 321326 106634
rect 321562 106398 321646 106634
rect 321882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 64826 102454
rect 65062 102218 65146 102454
rect 65382 102218 100826 102454
rect 101062 102218 101146 102454
rect 101382 102218 208826 102454
rect 209062 102218 209146 102454
rect 209382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 316826 102454
rect 317062 102218 317146 102454
rect 317382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 64826 102134
rect 65062 101898 65146 102134
rect 65382 101898 100826 102134
rect 101062 101898 101146 102134
rect 101382 101898 208826 102134
rect 209062 101898 209146 102134
rect 209382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 316826 102134
rect 317062 101898 317146 102134
rect 317382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 60326 97954
rect 60562 97718 60646 97954
rect 60882 97718 96326 97954
rect 96562 97718 96646 97954
rect 96882 97718 204326 97954
rect 204562 97718 204646 97954
rect 204882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 312326 97954
rect 312562 97718 312646 97954
rect 312882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 60326 97634
rect 60562 97398 60646 97634
rect 60882 97398 96326 97634
rect 96562 97398 96646 97634
rect 96882 97398 204326 97634
rect 204562 97398 204646 97634
rect 204882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 312326 97634
rect 312562 97398 312646 97634
rect 312882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 87326 88954
rect 87562 88718 87646 88954
rect 87882 88718 195326 88954
rect 195562 88718 195646 88954
rect 195882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 303326 88954
rect 303562 88718 303646 88954
rect 303882 88718 339326 88954
rect 339562 88718 339646 88954
rect 339882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 87326 88634
rect 87562 88398 87646 88634
rect 87882 88398 195326 88634
rect 195562 88398 195646 88634
rect 195882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 303326 88634
rect 303562 88398 303646 88634
rect 303882 88398 339326 88634
rect 339562 88398 339646 88634
rect 339882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 82826 84454
rect 83062 84218 83146 84454
rect 83382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 298826 84454
rect 299062 84218 299146 84454
rect 299382 84218 334826 84454
rect 335062 84218 335146 84454
rect 335382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 82826 84134
rect 83062 83898 83146 84134
rect 83382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 298826 84134
rect 299062 83898 299146 84134
rect 299382 83898 334826 84134
rect 335062 83898 335146 84134
rect 335382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 78326 79954
rect 78562 79718 78646 79954
rect 78882 79718 114326 79954
rect 114562 79718 114646 79954
rect 114882 79718 222326 79954
rect 222562 79718 222646 79954
rect 222882 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 330326 79954
rect 330562 79718 330646 79954
rect 330882 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 78326 79634
rect 78562 79398 78646 79634
rect 78882 79398 114326 79634
rect 114562 79398 114646 79634
rect 114882 79398 222326 79634
rect 222562 79398 222646 79634
rect 222882 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 330326 79634
rect 330562 79398 330646 79634
rect 330882 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 69326 70954
rect 69562 70718 69646 70954
rect 69882 70718 105326 70954
rect 105562 70718 105646 70954
rect 105882 70718 141326 70954
rect 141562 70718 141646 70954
rect 141882 70718 177326 70954
rect 177562 70718 177646 70954
rect 177882 70718 213326 70954
rect 213562 70718 213646 70954
rect 213882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 321326 70954
rect 321562 70718 321646 70954
rect 321882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 69326 70634
rect 69562 70398 69646 70634
rect 69882 70398 105326 70634
rect 105562 70398 105646 70634
rect 105882 70398 141326 70634
rect 141562 70398 141646 70634
rect 141882 70398 177326 70634
rect 177562 70398 177646 70634
rect 177882 70398 213326 70634
rect 213562 70398 213646 70634
rect 213882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 321326 70634
rect 321562 70398 321646 70634
rect 321882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 64826 66454
rect 65062 66218 65146 66454
rect 65382 66218 100826 66454
rect 101062 66218 101146 66454
rect 101382 66218 136826 66454
rect 137062 66218 137146 66454
rect 137382 66218 172826 66454
rect 173062 66218 173146 66454
rect 173382 66218 208826 66454
rect 209062 66218 209146 66454
rect 209382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 316826 66454
rect 317062 66218 317146 66454
rect 317382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 64826 66134
rect 65062 65898 65146 66134
rect 65382 65898 100826 66134
rect 101062 65898 101146 66134
rect 101382 65898 136826 66134
rect 137062 65898 137146 66134
rect 137382 65898 172826 66134
rect 173062 65898 173146 66134
rect 173382 65898 208826 66134
rect 209062 65898 209146 66134
rect 209382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 316826 66134
rect 317062 65898 317146 66134
rect 317382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 60326 61954
rect 60562 61718 60646 61954
rect 60882 61718 96326 61954
rect 96562 61718 96646 61954
rect 96882 61718 132326 61954
rect 132562 61718 132646 61954
rect 132882 61718 168326 61954
rect 168562 61718 168646 61954
rect 168882 61718 204326 61954
rect 204562 61718 204646 61954
rect 204882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 312326 61954
rect 312562 61718 312646 61954
rect 312882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 60326 61634
rect 60562 61398 60646 61634
rect 60882 61398 96326 61634
rect 96562 61398 96646 61634
rect 96882 61398 132326 61634
rect 132562 61398 132646 61634
rect 132882 61398 168326 61634
rect 168562 61398 168646 61634
rect 168882 61398 204326 61634
rect 204562 61398 204646 61634
rect 204882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 312326 61634
rect 312562 61398 312646 61634
rect 312882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use rlbp_macro  rlbp_macro0
timestamp 0
transform 1 0 120000 0 1 80000
box 0 0 70000 60000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 142000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 78000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 142000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 142000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 142000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 78000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 142000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 142000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 78000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 142000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 142000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 78000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 142000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 142000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 78000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 142000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 142000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 78000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 142000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 142000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 78000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 142000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 142000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 78000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 142000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
