magic
tech sky130A
magscale 1 2
timestamp 1668356327
<< nwell >>
rect 285 -700 1125 -375
<< pwell >>
rect 320 -785 1125 -780
rect 285 -975 1125 -785
<< nmos >>
rect 430 -910 460 -805
rect 535 -910 565 -805
rect 765 -910 795 -805
rect 995 -910 1025 -805
<< pmos >>
rect 430 -615 460 -460
rect 535 -615 565 -460
rect 760 -615 790 -460
rect 990 -615 1020 -460
<< ndiff >>
rect 365 -850 430 -805
rect 365 -885 380 -850
rect 415 -885 430 -850
rect 365 -910 430 -885
rect 460 -910 535 -805
rect 565 -845 625 -805
rect 565 -880 580 -845
rect 615 -880 625 -845
rect 565 -910 625 -880
rect 700 -850 765 -805
rect 700 -885 715 -850
rect 750 -885 765 -850
rect 700 -910 765 -885
rect 795 -845 855 -805
rect 795 -880 810 -845
rect 845 -880 855 -845
rect 795 -910 855 -880
rect 930 -850 995 -805
rect 930 -885 945 -850
rect 980 -885 995 -850
rect 930 -910 995 -885
rect 1025 -845 1085 -805
rect 1025 -880 1040 -845
rect 1075 -880 1085 -845
rect 1025 -910 1085 -880
<< pdiff >>
rect 370 -480 430 -460
rect 370 -515 380 -480
rect 415 -515 430 -480
rect 370 -550 430 -515
rect 370 -585 380 -550
rect 415 -585 430 -550
rect 370 -615 430 -585
rect 460 -615 535 -460
rect 565 -485 625 -460
rect 565 -520 580 -485
rect 615 -520 625 -485
rect 565 -560 625 -520
rect 565 -595 580 -560
rect 615 -595 625 -560
rect 565 -615 625 -595
rect 700 -480 760 -460
rect 700 -515 710 -480
rect 745 -515 760 -480
rect 700 -550 760 -515
rect 700 -585 710 -550
rect 745 -585 760 -550
rect 700 -615 760 -585
rect 790 -485 850 -460
rect 790 -520 805 -485
rect 840 -520 850 -485
rect 790 -560 850 -520
rect 790 -595 805 -560
rect 840 -595 850 -560
rect 790 -615 850 -595
rect 930 -480 990 -460
rect 930 -515 940 -480
rect 975 -515 990 -480
rect 930 -550 990 -515
rect 930 -585 940 -550
rect 975 -585 990 -550
rect 930 -615 990 -585
rect 1020 -485 1080 -460
rect 1020 -520 1035 -485
rect 1070 -520 1080 -485
rect 1020 -560 1080 -520
rect 1020 -595 1035 -560
rect 1070 -595 1080 -560
rect 1020 -615 1080 -595
<< ndiffc >>
rect 380 -885 415 -850
rect 580 -880 615 -845
rect 715 -885 750 -850
rect 810 -880 845 -845
rect 945 -885 980 -850
rect 1040 -880 1075 -845
<< pdiffc >>
rect 380 -515 415 -480
rect 380 -585 415 -550
rect 580 -520 615 -485
rect 580 -595 615 -560
rect 710 -515 745 -480
rect 710 -585 745 -550
rect 805 -520 840 -485
rect 805 -595 840 -560
rect 940 -515 975 -480
rect 940 -585 975 -550
rect 1035 -520 1070 -485
rect 1035 -595 1070 -560
<< poly >>
rect 430 -460 460 -430
rect 535 -460 565 -430
rect 760 -460 790 -430
rect 990 -460 1020 -430
rect 430 -650 460 -615
rect 400 -665 475 -650
rect 400 -700 420 -665
rect 455 -700 475 -665
rect 535 -700 565 -615
rect 760 -645 790 -615
rect 990 -645 1020 -615
rect 760 -665 795 -645
rect 990 -665 1025 -645
rect 740 -685 795 -665
rect 400 -710 475 -700
rect 520 -720 575 -700
rect 285 -735 360 -725
rect 285 -770 305 -735
rect 340 -755 360 -735
rect 520 -755 530 -720
rect 565 -755 575 -720
rect 740 -720 750 -685
rect 785 -720 795 -685
rect 740 -740 795 -720
rect 970 -685 1025 -665
rect 970 -720 980 -685
rect 1015 -720 1025 -685
rect 970 -740 1025 -720
rect 340 -770 460 -755
rect 285 -785 460 -770
rect 520 -775 575 -755
rect 760 -760 795 -740
rect 990 -760 1025 -740
rect 430 -805 460 -785
rect 535 -805 565 -775
rect 765 -805 795 -760
rect 995 -805 1025 -760
rect 430 -940 460 -910
rect 535 -940 565 -910
rect 765 -940 795 -910
rect 995 -940 1025 -910
<< polycont >>
rect 420 -700 455 -665
rect 305 -770 340 -735
rect 530 -755 565 -720
rect 750 -720 785 -685
rect 980 -720 1015 -685
<< locali >>
rect 285 -430 330 -395
rect 365 -430 425 -395
rect 460 -430 520 -395
rect 555 -430 615 -395
rect 650 -430 710 -395
rect 745 -430 805 -395
rect 840 -430 900 -395
rect 935 -430 995 -395
rect 1030 -430 1125 -395
rect 370 -480 425 -430
rect 370 -515 380 -480
rect 415 -515 425 -480
rect 370 -550 425 -515
rect 370 -585 380 -550
rect 415 -585 425 -550
rect 370 -610 425 -585
rect 570 -485 625 -465
rect 570 -520 580 -485
rect 615 -520 625 -485
rect 570 -560 625 -520
rect 570 -595 580 -560
rect 615 -595 625 -560
rect 570 -615 625 -595
rect 700 -480 755 -430
rect 700 -515 710 -480
rect 745 -515 755 -480
rect 700 -550 755 -515
rect 700 -585 710 -550
rect 745 -585 755 -550
rect 700 -615 755 -585
rect 795 -470 850 -465
rect 795 -485 870 -470
rect 795 -520 805 -485
rect 840 -520 870 -485
rect 795 -560 870 -520
rect 795 -595 805 -560
rect 840 -595 870 -560
rect 795 -615 870 -595
rect 930 -480 985 -430
rect 930 -515 940 -480
rect 975 -515 985 -480
rect 930 -550 985 -515
rect 930 -585 940 -550
rect 975 -585 985 -550
rect 930 -615 985 -585
rect 1025 -470 1080 -465
rect 1025 -485 1100 -470
rect 1025 -520 1035 -485
rect 1070 -520 1100 -485
rect 1025 -560 1100 -520
rect 1025 -595 1035 -560
rect 1070 -595 1100 -560
rect 1025 -615 1100 -595
rect 400 -665 475 -650
rect 570 -655 655 -615
rect 400 -700 415 -665
rect 455 -700 475 -665
rect 620 -690 655 -655
rect 740 -685 795 -665
rect 740 -690 750 -685
rect 400 -710 475 -700
rect 520 -720 575 -700
rect 285 -735 360 -725
rect 285 -770 305 -735
rect 340 -770 360 -735
rect 285 -785 360 -770
rect 520 -755 530 -720
rect 565 -755 575 -720
rect 520 -775 575 -755
rect 620 -720 750 -690
rect 785 -720 795 -685
rect 620 -735 795 -720
rect 620 -810 655 -735
rect 740 -740 795 -735
rect 835 -700 870 -615
rect 970 -685 1025 -665
rect 970 -700 980 -685
rect 835 -720 980 -700
rect 1015 -720 1025 -685
rect 835 -740 1025 -720
rect 835 -780 870 -740
rect 1065 -775 1100 -615
rect 375 -850 420 -820
rect 375 -885 380 -850
rect 415 -885 420 -850
rect 375 -940 420 -885
rect 570 -845 655 -810
rect 805 -820 870 -780
rect 1035 -785 1110 -775
rect 1035 -820 1055 -785
rect 1090 -820 1110 -785
rect 570 -880 580 -845
rect 615 -855 655 -845
rect 710 -850 755 -820
rect 615 -880 630 -855
rect 570 -900 630 -880
rect 710 -885 715 -850
rect 750 -885 755 -850
rect 710 -940 755 -885
rect 805 -845 850 -820
rect 805 -880 810 -845
rect 845 -880 850 -845
rect 805 -900 850 -880
rect 940 -850 985 -820
rect 940 -885 945 -850
rect 980 -885 985 -850
rect 940 -940 985 -885
rect 1035 -830 1110 -820
rect 1035 -845 1080 -830
rect 1035 -880 1040 -845
rect 1075 -880 1080 -845
rect 1035 -900 1080 -880
rect 285 -975 330 -940
rect 365 -975 425 -940
rect 460 -975 520 -940
rect 555 -975 615 -940
rect 650 -975 710 -940
rect 745 -975 805 -940
rect 840 -975 900 -940
rect 935 -975 995 -940
rect 1030 -975 1125 -940
<< viali >>
rect 330 -430 365 -395
rect 425 -430 460 -395
rect 520 -430 555 -395
rect 615 -430 650 -395
rect 710 -430 745 -395
rect 805 -430 840 -395
rect 900 -430 935 -395
rect 995 -430 1030 -395
rect 415 -700 420 -665
rect 420 -700 455 -665
rect 530 -755 565 -720
rect 750 -720 785 -685
rect 1055 -820 1090 -785
rect 330 -975 365 -940
rect 425 -975 460 -940
rect 520 -975 555 -940
rect 615 -975 650 -940
rect 710 -975 745 -940
rect 805 -975 840 -940
rect 900 -975 935 -940
rect 995 -975 1030 -940
<< metal1 >>
rect 304 397 499 403
rect 304 -200 499 202
rect 300 -365 500 -200
rect 275 -395 1125 -365
rect 275 -430 330 -395
rect 365 -430 425 -395
rect 460 -430 520 -395
rect 555 -430 615 -395
rect 650 -430 710 -395
rect 745 -430 805 -395
rect 840 -430 900 -395
rect 935 -430 995 -395
rect 1030 -430 1125 -395
rect 275 -460 1125 -430
rect -540 -545 -120 -490
rect -540 -595 345 -545
rect -540 -650 -120 -595
rect 295 -610 345 -595
rect 295 -650 450 -610
rect 295 -660 475 -650
rect 400 -665 475 -660
rect -540 -730 -120 -690
rect 400 -700 415 -665
rect 455 -700 475 -665
rect 740 -685 795 -665
rect 400 -710 475 -700
rect 520 -720 575 -700
rect 285 -730 360 -725
rect -540 -780 360 -730
rect -540 -850 -120 -780
rect 285 -785 360 -780
rect 520 -755 530 -720
rect 565 -740 575 -720
rect 740 -720 750 -685
rect 785 -705 795 -685
rect 785 -720 850 -705
rect 740 -740 850 -720
rect 565 -755 580 -740
rect 520 -800 580 -755
rect 820 -790 850 -740
rect 1035 -785 1110 -775
rect 1035 -790 1055 -785
rect 520 -827 565 -800
rect 820 -820 1055 -790
rect 1090 -790 1110 -785
rect 1220 -790 1640 -720
rect 1090 -820 1640 -790
rect 8 -872 565 -827
rect 1035 -830 1110 -820
rect -540 -1067 -120 -1010
rect 8 -1067 53 -872
rect 1220 -880 1640 -820
rect 285 -940 1125 -910
rect 285 -975 330 -940
rect 365 -975 425 -940
rect 460 -975 520 -940
rect 555 -975 615 -940
rect 650 -975 710 -940
rect 745 -975 805 -940
rect 840 -975 900 -940
rect 935 -975 995 -940
rect 1030 -975 1125 -940
rect 285 -1005 1125 -975
rect -540 -1112 53 -1067
rect -540 -1170 -120 -1112
rect 300 -1500 500 -1005
rect 300 -1706 500 -1700
<< via1 >>
rect 304 202 499 397
rect 300 -1700 500 -1500
<< metal2 >>
rect 200 397 600 500
rect 200 202 304 397
rect 499 202 600 397
rect 200 100 600 202
rect 200 -1500 600 -1400
rect 200 -1700 300 -1500
rect 500 -1700 600 -1500
rect 200 -1800 600 -1700
<< via2 >>
rect 304 202 499 397
rect 300 -1700 500 -1500
<< metal3 >>
rect 200 402 600 500
rect 200 197 299 402
rect 504 197 600 402
rect 200 100 600 197
rect 200 -1495 600 -1400
rect 200 -1705 295 -1495
rect 505 -1705 600 -1495
rect 200 -1800 600 -1705
<< via3 >>
rect 299 397 504 402
rect 299 202 304 397
rect 304 202 499 397
rect 499 202 504 397
rect 299 197 504 202
rect 295 -1500 505 -1495
rect 295 -1700 300 -1500
rect 300 -1700 500 -1500
rect 500 -1700 505 -1500
rect 295 -1705 505 -1700
<< metal4 >>
rect -100 900 2200 1600
rect 304 403 499 900
rect 298 402 505 403
rect 298 197 299 402
rect 504 197 505 402
rect 298 196 505 197
rect 294 -1495 506 -1494
rect 294 -1705 295 -1495
rect 505 -1705 506 -1495
rect 294 -1706 506 -1705
rect 300 -2200 500 -1706
rect -100 -2900 2200 -2200
<< labels >>
flabel metal1 285 -960 285 -960 0 FreeSans 80 0 0 0 VSS
port 0 nsew ground input
flabel metal1 275 -415 275 -415 0 FreeSans 80 0 0 0 VDD
port 1 nsew power input
flabel metal1 405 -685 405 -685 0 FreeSans 80 0 0 0 M
port 2 nsew signal input
flabel metal1 290 -760 290 -760 0 FreeSans 80 0 0 0 P
port 3 nsew signal input
flabel metal1 525 -740 525 -740 0 FreeSans 80 0 0 0 C
port 4 nsew signal input
flabel metal1 1105 -805 1105 -805 0 FreeSans 80 0 0 0 OUT
port 5 nsew signal output
<< end >>
